
module pipeline ( clock, reset, fake_out );
  input clock, reset;
  output fake_out;
  wire   stall, wrenable, jal_0, mem2reg_1, regwrite_1, jal_1, regwrite_2,
         jal_2, stallack, N14, N15, N17, N19, N23, N27, N28, N32, N34, N38,
         N43, N44, N46, N47, N139, decode_N4, decode_N2, decode_rs2_0_,
         decode_rs2_1_, decode_rs2_2_, decode_rs2_3_, decode_rs2_4_,
         decode_rs1_2_, decode_rs1_3_, decode_rs1_4_, decode_decoder_N279,
         decode_decoder_N278, decode_decoder_N277, decode_decoder_N276,
         decode_decoder_N275, decode_decoder_N274, decode_decoder_N273,
         decode_regfile_N163, decode_regfile_N162, decode_regfile_N161,
         decode_regfile_N160, decode_regfile_N159, decode_regfile_N158,
         decode_regfile_N157, decode_regfile_N156, decode_regfile_N155,
         decode_regfile_N154, decode_regfile_N153, decode_regfile_N152,
         decode_regfile_N151, decode_regfile_N150, decode_regfile_N149,
         decode_regfile_N148, decode_regfile_N147, decode_regfile_N146,
         decode_regfile_N145, decode_regfile_N144, decode_regfile_N143,
         decode_regfile_N142, decode_regfile_N141, decode_regfile_N140,
         decode_regfile_N139, decode_regfile_N138, decode_regfile_N137,
         decode_regfile_N136, decode_regfile_N135, decode_regfile_N134,
         decode_regfile_N133, decode_regfile_N132, decode_regfile_N131,
         decode_regfile_N130, decode_regfile_N129, decode_regfile_N128,
         decode_regfile_N127, decode_regfile_N126, decode_regfile_N125,
         decode_regfile_N124, decode_regfile_N123, decode_regfile_N122,
         decode_regfile_N121, decode_regfile_N120, decode_regfile_N119,
         decode_regfile_N118, decode_regfile_N117, decode_regfile_N116,
         decode_regfile_N115, decode_regfile_N114, decode_regfile_N113,
         decode_regfile_N112, decode_regfile_N111, decode_regfile_N110,
         decode_regfile_N109, decode_regfile_N108, decode_regfile_N107,
         decode_regfile_N106, decode_regfile_N105, decode_regfile_N104,
         decode_regfile_N103, decode_regfile_N102, decode_regfile_N101,
         decode_regfile_N100, decode_regfile_N91, decode_regfile_N90,
         decode_regfile_N89, decode_regfile_N88, decode_regfile_N87,
         decode_regfile_N86, decode_regfile_N85, decode_regfile_N84,
         decode_regfile_N83, decode_regfile_N82, decode_regfile_N81,
         decode_regfile_N80, decode_regfile_N79, decode_regfile_N78,
         decode_regfile_N77, decode_regfile_N76, decode_regfile_N75,
         decode_regfile_N74, decode_regfile_N73, decode_regfile_N72,
         decode_regfile_N71, decode_regfile_N70, decode_regfile_N69,
         decode_regfile_N68, decode_regfile_N67, decode_regfile_N66,
         decode_regfile_N65, decode_regfile_N64, decode_regfile_N63,
         decode_regfile_N62, decode_regfile_N61, decode_regfile_N60,
         decode_regfile_N59, decode_regfile_N58, decode_regfile_N57,
         decode_regfile_N56, decode_regfile_N55, decode_regfile_N54,
         decode_regfile_N53, decode_regfile_N52, decode_regfile_N51,
         decode_regfile_N50, decode_regfile_N49, decode_regfile_N48,
         decode_regfile_N47, decode_regfile_N46, decode_regfile_N45,
         decode_regfile_N44, decode_regfile_N43, decode_regfile_N42,
         decode_regfile_N41, decode_regfile_N40, decode_regfile_N39,
         decode_regfile_N38, decode_regfile_N37, decode_regfile_N36,
         decode_regfile_N35, decode_regfile_N34, decode_regfile_N33,
         decode_regfile_N32, decode_regfile_N31, decode_regfile_N30,
         decode_regfile_N29, decode_regfile_N28, decode_regfile_intregs_0__0_,
         decode_regfile_intregs_0__1_, decode_regfile_intregs_0__2_,
         decode_regfile_intregs_0__3_, decode_regfile_intregs_0__4_,
         decode_regfile_intregs_0__5_, decode_regfile_intregs_0__6_,
         decode_regfile_intregs_0__7_, decode_regfile_intregs_0__8_,
         decode_regfile_intregs_0__9_, decode_regfile_intregs_0__10_,
         decode_regfile_intregs_0__11_, decode_regfile_intregs_0__12_,
         decode_regfile_intregs_0__13_, decode_regfile_intregs_0__14_,
         decode_regfile_intregs_0__15_, decode_regfile_intregs_0__16_,
         decode_regfile_intregs_0__17_, decode_regfile_intregs_0__18_,
         decode_regfile_intregs_0__19_, decode_regfile_intregs_0__20_,
         decode_regfile_intregs_0__21_, decode_regfile_intregs_0__22_,
         decode_regfile_intregs_0__23_, decode_regfile_intregs_0__24_,
         decode_regfile_intregs_0__25_, decode_regfile_intregs_0__26_,
         decode_regfile_intregs_0__27_, decode_regfile_intregs_0__28_,
         decode_regfile_intregs_0__29_, decode_regfile_intregs_0__30_,
         decode_regfile_intregs_0__31_, decode_regfile_intregs_1__0_,
         decode_regfile_intregs_1__1_, decode_regfile_intregs_1__2_,
         decode_regfile_intregs_1__3_, decode_regfile_intregs_1__4_,
         decode_regfile_intregs_1__5_, decode_regfile_intregs_1__6_,
         decode_regfile_intregs_1__7_, decode_regfile_intregs_1__8_,
         decode_regfile_intregs_1__9_, decode_regfile_intregs_1__10_,
         decode_regfile_intregs_1__11_, decode_regfile_intregs_1__12_,
         decode_regfile_intregs_1__13_, decode_regfile_intregs_1__14_,
         decode_regfile_intregs_1__15_, decode_regfile_intregs_1__16_,
         decode_regfile_intregs_1__17_, decode_regfile_intregs_1__18_,
         decode_regfile_intregs_1__19_, decode_regfile_intregs_1__20_,
         decode_regfile_intregs_1__21_, decode_regfile_intregs_1__22_,
         decode_regfile_intregs_1__23_, decode_regfile_intregs_1__24_,
         decode_regfile_intregs_1__25_, decode_regfile_intregs_1__26_,
         decode_regfile_intregs_1__27_, decode_regfile_intregs_1__28_,
         decode_regfile_intregs_1__29_, decode_regfile_intregs_1__30_,
         decode_regfile_intregs_1__31_, decode_regfile_intregs_2__0_,
         decode_regfile_intregs_2__1_, decode_regfile_intregs_2__2_,
         decode_regfile_intregs_2__3_, decode_regfile_intregs_2__4_,
         decode_regfile_intregs_2__5_, decode_regfile_intregs_2__6_,
         decode_regfile_intregs_2__7_, decode_regfile_intregs_2__8_,
         decode_regfile_intregs_2__9_, decode_regfile_intregs_2__10_,
         decode_regfile_intregs_2__11_, decode_regfile_intregs_2__12_,
         decode_regfile_intregs_2__13_, decode_regfile_intregs_2__14_,
         decode_regfile_intregs_2__15_, decode_regfile_intregs_2__16_,
         decode_regfile_intregs_2__17_, decode_regfile_intregs_2__18_,
         decode_regfile_intregs_2__19_, decode_regfile_intregs_2__20_,
         decode_regfile_intregs_2__21_, decode_regfile_intregs_2__22_,
         decode_regfile_intregs_2__23_, decode_regfile_intregs_2__24_,
         decode_regfile_intregs_2__25_, decode_regfile_intregs_2__26_,
         decode_regfile_intregs_2__27_, decode_regfile_intregs_2__28_,
         decode_regfile_intregs_2__29_, decode_regfile_intregs_2__30_,
         decode_regfile_intregs_2__31_, decode_regfile_intregs_3__0_,
         decode_regfile_intregs_3__1_, decode_regfile_intregs_3__2_,
         decode_regfile_intregs_3__3_, decode_regfile_intregs_3__4_,
         decode_regfile_intregs_3__5_, decode_regfile_intregs_3__6_,
         decode_regfile_intregs_3__7_, decode_regfile_intregs_3__8_,
         decode_regfile_intregs_3__9_, decode_regfile_intregs_3__10_,
         decode_regfile_intregs_3__11_, decode_regfile_intregs_3__12_,
         decode_regfile_intregs_3__13_, decode_regfile_intregs_3__14_,
         decode_regfile_intregs_3__15_, decode_regfile_intregs_3__16_,
         decode_regfile_intregs_3__17_, decode_regfile_intregs_3__18_,
         decode_regfile_intregs_3__19_, decode_regfile_intregs_3__20_,
         decode_regfile_intregs_3__21_, decode_regfile_intregs_3__22_,
         decode_regfile_intregs_3__23_, decode_regfile_intregs_3__24_,
         decode_regfile_intregs_3__25_, decode_regfile_intregs_3__26_,
         decode_regfile_intregs_3__27_, decode_regfile_intregs_3__28_,
         decode_regfile_intregs_3__29_, decode_regfile_intregs_3__30_,
         decode_regfile_intregs_3__31_, decode_regfile_intregs_4__0_,
         decode_regfile_intregs_4__1_, decode_regfile_intregs_4__2_,
         decode_regfile_intregs_4__3_, decode_regfile_intregs_4__4_,
         decode_regfile_intregs_4__5_, decode_regfile_intregs_4__6_,
         decode_regfile_intregs_4__7_, decode_regfile_intregs_4__8_,
         decode_regfile_intregs_4__9_, decode_regfile_intregs_4__10_,
         decode_regfile_intregs_4__11_, decode_regfile_intregs_4__12_,
         decode_regfile_intregs_4__13_, decode_regfile_intregs_4__14_,
         decode_regfile_intregs_4__15_, decode_regfile_intregs_4__16_,
         decode_regfile_intregs_4__17_, decode_regfile_intregs_4__18_,
         decode_regfile_intregs_4__19_, decode_regfile_intregs_4__20_,
         decode_regfile_intregs_4__21_, decode_regfile_intregs_4__22_,
         decode_regfile_intregs_4__23_, decode_regfile_intregs_4__24_,
         decode_regfile_intregs_4__25_, decode_regfile_intregs_4__26_,
         decode_regfile_intregs_4__27_, decode_regfile_intregs_4__28_,
         decode_regfile_intregs_4__29_, decode_regfile_intregs_4__30_,
         decode_regfile_intregs_4__31_, decode_regfile_intregs_5__0_,
         decode_regfile_intregs_5__1_, decode_regfile_intregs_5__2_,
         decode_regfile_intregs_5__3_, decode_regfile_intregs_5__4_,
         decode_regfile_intregs_5__5_, decode_regfile_intregs_5__6_,
         decode_regfile_intregs_5__7_, decode_regfile_intregs_5__8_,
         decode_regfile_intregs_5__9_, decode_regfile_intregs_5__10_,
         decode_regfile_intregs_5__11_, decode_regfile_intregs_5__12_,
         decode_regfile_intregs_5__13_, decode_regfile_intregs_5__14_,
         decode_regfile_intregs_5__15_, decode_regfile_intregs_5__16_,
         decode_regfile_intregs_5__17_, decode_regfile_intregs_5__18_,
         decode_regfile_intregs_5__19_, decode_regfile_intregs_5__20_,
         decode_regfile_intregs_5__21_, decode_regfile_intregs_5__22_,
         decode_regfile_intregs_5__23_, decode_regfile_intregs_5__24_,
         decode_regfile_intregs_5__25_, decode_regfile_intregs_5__26_,
         decode_regfile_intregs_5__27_, decode_regfile_intregs_5__28_,
         decode_regfile_intregs_5__29_, decode_regfile_intregs_5__30_,
         decode_regfile_intregs_5__31_, decode_regfile_intregs_6__0_,
         decode_regfile_intregs_6__1_, decode_regfile_intregs_6__2_,
         decode_regfile_intregs_6__3_, decode_regfile_intregs_6__4_,
         decode_regfile_intregs_6__5_, decode_regfile_intregs_6__6_,
         decode_regfile_intregs_6__7_, decode_regfile_intregs_6__8_,
         decode_regfile_intregs_6__9_, decode_regfile_intregs_6__10_,
         decode_regfile_intregs_6__11_, decode_regfile_intregs_6__12_,
         decode_regfile_intregs_6__13_, decode_regfile_intregs_6__14_,
         decode_regfile_intregs_6__15_, decode_regfile_intregs_6__16_,
         decode_regfile_intregs_6__17_, decode_regfile_intregs_6__18_,
         decode_regfile_intregs_6__19_, decode_regfile_intregs_6__20_,
         decode_regfile_intregs_6__21_, decode_regfile_intregs_6__22_,
         decode_regfile_intregs_6__23_, decode_regfile_intregs_6__24_,
         decode_regfile_intregs_6__25_, decode_regfile_intregs_6__26_,
         decode_regfile_intregs_6__27_, decode_regfile_intregs_6__28_,
         decode_regfile_intregs_6__29_, decode_regfile_intregs_6__30_,
         decode_regfile_intregs_6__31_, decode_regfile_intregs_7__0_,
         decode_regfile_intregs_7__1_, decode_regfile_intregs_7__2_,
         decode_regfile_intregs_7__3_, decode_regfile_intregs_7__4_,
         decode_regfile_intregs_7__5_, decode_regfile_intregs_7__6_,
         decode_regfile_intregs_7__7_, decode_regfile_intregs_7__8_,
         decode_regfile_intregs_7__9_, decode_regfile_intregs_7__10_,
         decode_regfile_intregs_7__11_, decode_regfile_intregs_7__12_,
         decode_regfile_intregs_7__13_, decode_regfile_intregs_7__14_,
         decode_regfile_intregs_7__15_, decode_regfile_intregs_7__16_,
         decode_regfile_intregs_7__17_, decode_regfile_intregs_7__18_,
         decode_regfile_intregs_7__19_, decode_regfile_intregs_7__20_,
         decode_regfile_intregs_7__21_, decode_regfile_intregs_7__22_,
         decode_regfile_intregs_7__23_, decode_regfile_intregs_7__24_,
         decode_regfile_intregs_7__25_, decode_regfile_intregs_7__26_,
         decode_regfile_intregs_7__27_, decode_regfile_intregs_7__28_,
         decode_regfile_intregs_7__29_, decode_regfile_intregs_7__30_,
         decode_regfile_intregs_7__31_, decode_regfile_intregs_8__0_,
         decode_regfile_intregs_8__1_, decode_regfile_intregs_8__2_,
         decode_regfile_intregs_8__3_, decode_regfile_intregs_8__4_,
         decode_regfile_intregs_8__5_, decode_regfile_intregs_8__6_,
         decode_regfile_intregs_8__7_, decode_regfile_intregs_8__8_,
         decode_regfile_intregs_8__9_, decode_regfile_intregs_8__10_,
         decode_regfile_intregs_8__11_, decode_regfile_intregs_8__12_,
         decode_regfile_intregs_8__13_, decode_regfile_intregs_8__14_,
         decode_regfile_intregs_8__15_, decode_regfile_intregs_8__16_,
         decode_regfile_intregs_8__17_, decode_regfile_intregs_8__18_,
         decode_regfile_intregs_8__19_, decode_regfile_intregs_8__20_,
         decode_regfile_intregs_8__21_, decode_regfile_intregs_8__22_,
         decode_regfile_intregs_8__23_, decode_regfile_intregs_8__24_,
         decode_regfile_intregs_8__25_, decode_regfile_intregs_8__26_,
         decode_regfile_intregs_8__27_, decode_regfile_intregs_8__28_,
         decode_regfile_intregs_8__29_, decode_regfile_intregs_8__30_,
         decode_regfile_intregs_8__31_, decode_regfile_intregs_9__0_,
         decode_regfile_intregs_9__1_, decode_regfile_intregs_9__2_,
         decode_regfile_intregs_9__3_, decode_regfile_intregs_9__4_,
         decode_regfile_intregs_9__5_, decode_regfile_intregs_9__6_,
         decode_regfile_intregs_9__7_, decode_regfile_intregs_9__8_,
         decode_regfile_intregs_9__9_, decode_regfile_intregs_9__10_,
         decode_regfile_intregs_9__11_, decode_regfile_intregs_9__12_,
         decode_regfile_intregs_9__13_, decode_regfile_intregs_9__14_,
         decode_regfile_intregs_9__15_, decode_regfile_intregs_9__16_,
         decode_regfile_intregs_9__17_, decode_regfile_intregs_9__18_,
         decode_regfile_intregs_9__19_, decode_regfile_intregs_9__20_,
         decode_regfile_intregs_9__21_, decode_regfile_intregs_9__22_,
         decode_regfile_intregs_9__23_, decode_regfile_intregs_9__24_,
         decode_regfile_intregs_9__25_, decode_regfile_intregs_9__26_,
         decode_regfile_intregs_9__27_, decode_regfile_intregs_9__28_,
         decode_regfile_intregs_9__29_, decode_regfile_intregs_9__30_,
         decode_regfile_intregs_9__31_, decode_regfile_intregs_10__0_,
         decode_regfile_intregs_10__1_, decode_regfile_intregs_10__2_,
         decode_regfile_intregs_10__3_, decode_regfile_intregs_10__4_,
         decode_regfile_intregs_10__5_, decode_regfile_intregs_10__6_,
         decode_regfile_intregs_10__7_, decode_regfile_intregs_10__8_,
         decode_regfile_intregs_10__9_, decode_regfile_intregs_10__10_,
         decode_regfile_intregs_10__11_, decode_regfile_intregs_10__12_,
         decode_regfile_intregs_10__13_, decode_regfile_intregs_10__14_,
         decode_regfile_intregs_10__15_, decode_regfile_intregs_10__16_,
         decode_regfile_intregs_10__17_, decode_regfile_intregs_10__18_,
         decode_regfile_intregs_10__19_, decode_regfile_intregs_10__20_,
         decode_regfile_intregs_10__21_, decode_regfile_intregs_10__22_,
         decode_regfile_intregs_10__23_, decode_regfile_intregs_10__24_,
         decode_regfile_intregs_10__25_, decode_regfile_intregs_10__26_,
         decode_regfile_intregs_10__27_, decode_regfile_intregs_10__28_,
         decode_regfile_intregs_10__29_, decode_regfile_intregs_10__30_,
         decode_regfile_intregs_10__31_, decode_regfile_intregs_11__0_,
         decode_regfile_intregs_11__1_, decode_regfile_intregs_11__2_,
         decode_regfile_intregs_11__3_, decode_regfile_intregs_11__4_,
         decode_regfile_intregs_11__5_, decode_regfile_intregs_11__6_,
         decode_regfile_intregs_11__7_, decode_regfile_intregs_11__8_,
         decode_regfile_intregs_11__9_, decode_regfile_intregs_11__10_,
         decode_regfile_intregs_11__11_, decode_regfile_intregs_11__12_,
         decode_regfile_intregs_11__13_, decode_regfile_intregs_11__14_,
         decode_regfile_intregs_11__15_, decode_regfile_intregs_11__16_,
         decode_regfile_intregs_11__17_, decode_regfile_intregs_11__18_,
         decode_regfile_intregs_11__19_, decode_regfile_intregs_11__20_,
         decode_regfile_intregs_11__21_, decode_regfile_intregs_11__22_,
         decode_regfile_intregs_11__23_, decode_regfile_intregs_11__24_,
         decode_regfile_intregs_11__25_, decode_regfile_intregs_11__26_,
         decode_regfile_intregs_11__27_, decode_regfile_intregs_11__28_,
         decode_regfile_intregs_11__29_, decode_regfile_intregs_11__30_,
         decode_regfile_intregs_11__31_, decode_regfile_intregs_12__0_,
         decode_regfile_intregs_12__1_, decode_regfile_intregs_12__2_,
         decode_regfile_intregs_12__3_, decode_regfile_intregs_12__4_,
         decode_regfile_intregs_12__5_, decode_regfile_intregs_12__6_,
         decode_regfile_intregs_12__7_, decode_regfile_intregs_12__8_,
         decode_regfile_intregs_12__9_, decode_regfile_intregs_12__10_,
         decode_regfile_intregs_12__11_, decode_regfile_intregs_12__12_,
         decode_regfile_intregs_12__13_, decode_regfile_intregs_12__14_,
         decode_regfile_intregs_12__15_, decode_regfile_intregs_12__16_,
         decode_regfile_intregs_12__17_, decode_regfile_intregs_12__18_,
         decode_regfile_intregs_12__19_, decode_regfile_intregs_12__20_,
         decode_regfile_intregs_12__21_, decode_regfile_intregs_12__22_,
         decode_regfile_intregs_12__23_, decode_regfile_intregs_12__24_,
         decode_regfile_intregs_12__25_, decode_regfile_intregs_12__26_,
         decode_regfile_intregs_12__27_, decode_regfile_intregs_12__28_,
         decode_regfile_intregs_12__29_, decode_regfile_intregs_12__30_,
         decode_regfile_intregs_12__31_, decode_regfile_intregs_13__0_,
         decode_regfile_intregs_13__1_, decode_regfile_intregs_13__2_,
         decode_regfile_intregs_13__3_, decode_regfile_intregs_13__4_,
         decode_regfile_intregs_13__5_, decode_regfile_intregs_13__6_,
         decode_regfile_intregs_13__7_, decode_regfile_intregs_13__8_,
         decode_regfile_intregs_13__9_, decode_regfile_intregs_13__10_,
         decode_regfile_intregs_13__11_, decode_regfile_intregs_13__12_,
         decode_regfile_intregs_13__13_, decode_regfile_intregs_13__14_,
         decode_regfile_intregs_13__15_, decode_regfile_intregs_13__16_,
         decode_regfile_intregs_13__17_, decode_regfile_intregs_13__18_,
         decode_regfile_intregs_13__19_, decode_regfile_intregs_13__20_,
         decode_regfile_intregs_13__21_, decode_regfile_intregs_13__22_,
         decode_regfile_intregs_13__23_, decode_regfile_intregs_13__24_,
         decode_regfile_intregs_13__25_, decode_regfile_intregs_13__26_,
         decode_regfile_intregs_13__27_, decode_regfile_intregs_13__28_,
         decode_regfile_intregs_13__29_, decode_regfile_intregs_13__30_,
         decode_regfile_intregs_13__31_, decode_regfile_intregs_14__0_,
         decode_regfile_intregs_14__1_, decode_regfile_intregs_14__2_,
         decode_regfile_intregs_14__3_, decode_regfile_intregs_14__4_,
         decode_regfile_intregs_14__5_, decode_regfile_intregs_14__6_,
         decode_regfile_intregs_14__7_, decode_regfile_intregs_14__8_,
         decode_regfile_intregs_14__9_, decode_regfile_intregs_14__10_,
         decode_regfile_intregs_14__11_, decode_regfile_intregs_14__12_,
         decode_regfile_intregs_14__13_, decode_regfile_intregs_14__14_,
         decode_regfile_intregs_14__15_, decode_regfile_intregs_14__16_,
         decode_regfile_intregs_14__17_, decode_regfile_intregs_14__18_,
         decode_regfile_intregs_14__19_, decode_regfile_intregs_14__20_,
         decode_regfile_intregs_14__21_, decode_regfile_intregs_14__22_,
         decode_regfile_intregs_14__23_, decode_regfile_intregs_14__24_,
         decode_regfile_intregs_14__25_, decode_regfile_intregs_14__26_,
         decode_regfile_intregs_14__27_, decode_regfile_intregs_14__28_,
         decode_regfile_intregs_14__29_, decode_regfile_intregs_14__30_,
         decode_regfile_intregs_14__31_, decode_regfile_intregs_15__0_,
         decode_regfile_intregs_15__1_, decode_regfile_intregs_15__2_,
         decode_regfile_intregs_15__3_, decode_regfile_intregs_15__4_,
         decode_regfile_intregs_15__5_, decode_regfile_intregs_15__6_,
         decode_regfile_intregs_15__7_, decode_regfile_intregs_15__8_,
         decode_regfile_intregs_15__9_, decode_regfile_intregs_15__10_,
         decode_regfile_intregs_15__11_, decode_regfile_intregs_15__12_,
         decode_regfile_intregs_15__13_, decode_regfile_intregs_15__14_,
         decode_regfile_intregs_15__15_, decode_regfile_intregs_15__16_,
         decode_regfile_intregs_15__17_, decode_regfile_intregs_15__18_,
         decode_regfile_intregs_15__19_, decode_regfile_intregs_15__20_,
         decode_regfile_intregs_15__21_, decode_regfile_intregs_15__22_,
         decode_regfile_intregs_15__23_, decode_regfile_intregs_15__24_,
         decode_regfile_intregs_15__25_, decode_regfile_intregs_15__26_,
         decode_regfile_intregs_15__27_, decode_regfile_intregs_15__28_,
         decode_regfile_intregs_15__29_, decode_regfile_intregs_15__30_,
         decode_regfile_intregs_15__31_, decode_regfile_intregs_16__0_,
         decode_regfile_intregs_16__1_, decode_regfile_intregs_16__2_,
         decode_regfile_intregs_16__3_, decode_regfile_intregs_16__4_,
         decode_regfile_intregs_16__5_, decode_regfile_intregs_16__6_,
         decode_regfile_intregs_16__7_, decode_regfile_intregs_16__8_,
         decode_regfile_intregs_16__9_, decode_regfile_intregs_16__10_,
         decode_regfile_intregs_16__11_, decode_regfile_intregs_16__12_,
         decode_regfile_intregs_16__13_, decode_regfile_intregs_16__14_,
         decode_regfile_intregs_16__15_, decode_regfile_intregs_16__16_,
         decode_regfile_intregs_16__17_, decode_regfile_intregs_16__18_,
         decode_regfile_intregs_16__19_, decode_regfile_intregs_16__20_,
         decode_regfile_intregs_16__21_, decode_regfile_intregs_16__22_,
         decode_regfile_intregs_16__23_, decode_regfile_intregs_16__24_,
         decode_regfile_intregs_16__25_, decode_regfile_intregs_16__26_,
         decode_regfile_intregs_16__27_, decode_regfile_intregs_16__28_,
         decode_regfile_intregs_16__29_, decode_regfile_intregs_16__30_,
         decode_regfile_intregs_16__31_, decode_regfile_intregs_17__0_,
         decode_regfile_intregs_17__1_, decode_regfile_intregs_17__2_,
         decode_regfile_intregs_17__3_, decode_regfile_intregs_17__4_,
         decode_regfile_intregs_17__5_, decode_regfile_intregs_17__6_,
         decode_regfile_intregs_17__7_, decode_regfile_intregs_17__8_,
         decode_regfile_intregs_17__9_, decode_regfile_intregs_17__10_,
         decode_regfile_intregs_17__11_, decode_regfile_intregs_17__12_,
         decode_regfile_intregs_17__13_, decode_regfile_intregs_17__14_,
         decode_regfile_intregs_17__15_, decode_regfile_intregs_17__16_,
         decode_regfile_intregs_17__17_, decode_regfile_intregs_17__18_,
         decode_regfile_intregs_17__19_, decode_regfile_intregs_17__20_,
         decode_regfile_intregs_17__21_, decode_regfile_intregs_17__22_,
         decode_regfile_intregs_17__23_, decode_regfile_intregs_17__24_,
         decode_regfile_intregs_17__25_, decode_regfile_intregs_17__26_,
         decode_regfile_intregs_17__27_, decode_regfile_intregs_17__28_,
         decode_regfile_intregs_17__29_, decode_regfile_intregs_17__30_,
         decode_regfile_intregs_17__31_, decode_regfile_intregs_18__0_,
         decode_regfile_intregs_18__1_, decode_regfile_intregs_18__2_,
         decode_regfile_intregs_18__3_, decode_regfile_intregs_18__4_,
         decode_regfile_intregs_18__5_, decode_regfile_intregs_18__6_,
         decode_regfile_intregs_18__7_, decode_regfile_intregs_18__8_,
         decode_regfile_intregs_18__9_, decode_regfile_intregs_18__10_,
         decode_regfile_intregs_18__11_, decode_regfile_intregs_18__12_,
         decode_regfile_intregs_18__13_, decode_regfile_intregs_18__14_,
         decode_regfile_intregs_18__15_, decode_regfile_intregs_18__16_,
         decode_regfile_intregs_18__17_, decode_regfile_intregs_18__18_,
         decode_regfile_intregs_18__19_, decode_regfile_intregs_18__20_,
         decode_regfile_intregs_18__21_, decode_regfile_intregs_18__22_,
         decode_regfile_intregs_18__23_, decode_regfile_intregs_18__24_,
         decode_regfile_intregs_18__25_, decode_regfile_intregs_18__26_,
         decode_regfile_intregs_18__27_, decode_regfile_intregs_18__28_,
         decode_regfile_intregs_18__29_, decode_regfile_intregs_18__30_,
         decode_regfile_intregs_18__31_, decode_regfile_intregs_19__0_,
         decode_regfile_intregs_19__1_, decode_regfile_intregs_19__2_,
         decode_regfile_intregs_19__3_, decode_regfile_intregs_19__4_,
         decode_regfile_intregs_19__5_, decode_regfile_intregs_19__6_,
         decode_regfile_intregs_19__7_, decode_regfile_intregs_19__8_,
         decode_regfile_intregs_19__9_, decode_regfile_intregs_19__10_,
         decode_regfile_intregs_19__11_, decode_regfile_intregs_19__12_,
         decode_regfile_intregs_19__13_, decode_regfile_intregs_19__14_,
         decode_regfile_intregs_19__15_, decode_regfile_intregs_19__16_,
         decode_regfile_intregs_19__17_, decode_regfile_intregs_19__18_,
         decode_regfile_intregs_19__19_, decode_regfile_intregs_19__20_,
         decode_regfile_intregs_19__21_, decode_regfile_intregs_19__22_,
         decode_regfile_intregs_19__23_, decode_regfile_intregs_19__24_,
         decode_regfile_intregs_19__25_, decode_regfile_intregs_19__26_,
         decode_regfile_intregs_19__27_, decode_regfile_intregs_19__28_,
         decode_regfile_intregs_19__29_, decode_regfile_intregs_19__30_,
         decode_regfile_intregs_19__31_, decode_regfile_intregs_20__0_,
         decode_regfile_intregs_20__1_, decode_regfile_intregs_20__2_,
         decode_regfile_intregs_20__3_, decode_regfile_intregs_20__4_,
         decode_regfile_intregs_20__5_, decode_regfile_intregs_20__6_,
         decode_regfile_intregs_20__7_, decode_regfile_intregs_20__8_,
         decode_regfile_intregs_20__9_, decode_regfile_intregs_20__10_,
         decode_regfile_intregs_20__11_, decode_regfile_intregs_20__12_,
         decode_regfile_intregs_20__13_, decode_regfile_intregs_20__14_,
         decode_regfile_intregs_20__15_, decode_regfile_intregs_20__16_,
         decode_regfile_intregs_20__17_, decode_regfile_intregs_20__18_,
         decode_regfile_intregs_20__19_, decode_regfile_intregs_20__20_,
         decode_regfile_intregs_20__21_, decode_regfile_intregs_20__22_,
         decode_regfile_intregs_20__23_, decode_regfile_intregs_20__24_,
         decode_regfile_intregs_20__25_, decode_regfile_intregs_20__26_,
         decode_regfile_intregs_20__27_, decode_regfile_intregs_20__28_,
         decode_regfile_intregs_20__29_, decode_regfile_intregs_20__30_,
         decode_regfile_intregs_20__31_, decode_regfile_intregs_21__0_,
         decode_regfile_intregs_21__1_, decode_regfile_intregs_21__2_,
         decode_regfile_intregs_21__3_, decode_regfile_intregs_21__4_,
         decode_regfile_intregs_21__5_, decode_regfile_intregs_21__6_,
         decode_regfile_intregs_21__7_, decode_regfile_intregs_21__8_,
         decode_regfile_intregs_21__9_, decode_regfile_intregs_21__10_,
         decode_regfile_intregs_21__11_, decode_regfile_intregs_21__12_,
         decode_regfile_intregs_21__13_, decode_regfile_intregs_21__14_,
         decode_regfile_intregs_21__15_, decode_regfile_intregs_21__16_,
         decode_regfile_intregs_21__17_, decode_regfile_intregs_21__18_,
         decode_regfile_intregs_21__19_, decode_regfile_intregs_21__20_,
         decode_regfile_intregs_21__21_, decode_regfile_intregs_21__22_,
         decode_regfile_intregs_21__23_, decode_regfile_intregs_21__24_,
         decode_regfile_intregs_21__25_, decode_regfile_intregs_21__26_,
         decode_regfile_intregs_21__27_, decode_regfile_intregs_21__28_,
         decode_regfile_intregs_21__29_, decode_regfile_intregs_21__30_,
         decode_regfile_intregs_21__31_, decode_regfile_intregs_22__0_,
         decode_regfile_intregs_22__1_, decode_regfile_intregs_22__2_,
         decode_regfile_intregs_22__3_, decode_regfile_intregs_22__4_,
         decode_regfile_intregs_22__5_, decode_regfile_intregs_22__6_,
         decode_regfile_intregs_22__7_, decode_regfile_intregs_22__8_,
         decode_regfile_intregs_22__9_, decode_regfile_intregs_22__10_,
         decode_regfile_intregs_22__11_, decode_regfile_intregs_22__12_,
         decode_regfile_intregs_22__13_, decode_regfile_intregs_22__14_,
         decode_regfile_intregs_22__15_, decode_regfile_intregs_22__16_,
         decode_regfile_intregs_22__17_, decode_regfile_intregs_22__18_,
         decode_regfile_intregs_22__19_, decode_regfile_intregs_22__20_,
         decode_regfile_intregs_22__21_, decode_regfile_intregs_22__22_,
         decode_regfile_intregs_22__23_, decode_regfile_intregs_22__24_,
         decode_regfile_intregs_22__25_, decode_regfile_intregs_22__26_,
         decode_regfile_intregs_22__27_, decode_regfile_intregs_22__28_,
         decode_regfile_intregs_22__29_, decode_regfile_intregs_22__30_,
         decode_regfile_intregs_22__31_, decode_regfile_intregs_23__0_,
         decode_regfile_intregs_23__1_, decode_regfile_intregs_23__2_,
         decode_regfile_intregs_23__3_, decode_regfile_intregs_23__4_,
         decode_regfile_intregs_23__5_, decode_regfile_intregs_23__6_,
         decode_regfile_intregs_23__7_, decode_regfile_intregs_23__8_,
         decode_regfile_intregs_23__9_, decode_regfile_intregs_23__10_,
         decode_regfile_intregs_23__11_, decode_regfile_intregs_23__12_,
         decode_regfile_intregs_23__13_, decode_regfile_intregs_23__14_,
         decode_regfile_intregs_23__15_, decode_regfile_intregs_23__16_,
         decode_regfile_intregs_23__17_, decode_regfile_intregs_23__18_,
         decode_regfile_intregs_23__19_, decode_regfile_intregs_23__20_,
         decode_regfile_intregs_23__21_, decode_regfile_intregs_23__22_,
         decode_regfile_intregs_23__23_, decode_regfile_intregs_23__24_,
         decode_regfile_intregs_23__25_, decode_regfile_intregs_23__26_,
         decode_regfile_intregs_23__27_, decode_regfile_intregs_23__28_,
         decode_regfile_intregs_23__29_, decode_regfile_intregs_23__30_,
         decode_regfile_intregs_23__31_, decode_regfile_intregs_24__0_,
         decode_regfile_intregs_24__1_, decode_regfile_intregs_24__2_,
         decode_regfile_intregs_24__3_, decode_regfile_intregs_24__4_,
         decode_regfile_intregs_24__5_, decode_regfile_intregs_24__6_,
         decode_regfile_intregs_24__7_, decode_regfile_intregs_24__8_,
         decode_regfile_intregs_24__9_, decode_regfile_intregs_24__10_,
         decode_regfile_intregs_24__11_, decode_regfile_intregs_24__12_,
         decode_regfile_intregs_24__13_, decode_regfile_intregs_24__14_,
         decode_regfile_intregs_24__15_, decode_regfile_intregs_24__16_,
         decode_regfile_intregs_24__17_, decode_regfile_intregs_24__18_,
         decode_regfile_intregs_24__19_, decode_regfile_intregs_24__20_,
         decode_regfile_intregs_24__21_, decode_regfile_intregs_24__22_,
         decode_regfile_intregs_24__23_, decode_regfile_intregs_24__24_,
         decode_regfile_intregs_24__25_, decode_regfile_intregs_24__26_,
         decode_regfile_intregs_24__27_, decode_regfile_intregs_24__28_,
         decode_regfile_intregs_24__29_, decode_regfile_intregs_24__30_,
         decode_regfile_intregs_24__31_, decode_regfile_intregs_25__0_,
         decode_regfile_intregs_25__1_, decode_regfile_intregs_25__2_,
         decode_regfile_intregs_25__3_, decode_regfile_intregs_25__4_,
         decode_regfile_intregs_25__5_, decode_regfile_intregs_25__6_,
         decode_regfile_intregs_25__7_, decode_regfile_intregs_25__8_,
         decode_regfile_intregs_25__9_, decode_regfile_intregs_25__10_,
         decode_regfile_intregs_25__11_, decode_regfile_intregs_25__12_,
         decode_regfile_intregs_25__13_, decode_regfile_intregs_25__14_,
         decode_regfile_intregs_25__15_, decode_regfile_intregs_25__16_,
         decode_regfile_intregs_25__17_, decode_regfile_intregs_25__18_,
         decode_regfile_intregs_25__19_, decode_regfile_intregs_25__20_,
         decode_regfile_intregs_25__21_, decode_regfile_intregs_25__22_,
         decode_regfile_intregs_25__23_, decode_regfile_intregs_25__24_,
         decode_regfile_intregs_25__25_, decode_regfile_intregs_25__26_,
         decode_regfile_intregs_25__27_, decode_regfile_intregs_25__28_,
         decode_regfile_intregs_25__29_, decode_regfile_intregs_25__30_,
         decode_regfile_intregs_25__31_, decode_regfile_intregs_26__0_,
         decode_regfile_intregs_26__1_, decode_regfile_intregs_26__2_,
         decode_regfile_intregs_26__3_, decode_regfile_intregs_26__4_,
         decode_regfile_intregs_26__5_, decode_regfile_intregs_26__6_,
         decode_regfile_intregs_26__7_, decode_regfile_intregs_26__8_,
         decode_regfile_intregs_26__9_, decode_regfile_intregs_26__10_,
         decode_regfile_intregs_26__11_, decode_regfile_intregs_26__12_,
         decode_regfile_intregs_26__13_, decode_regfile_intregs_26__14_,
         decode_regfile_intregs_26__15_, decode_regfile_intregs_26__16_,
         decode_regfile_intregs_26__17_, decode_regfile_intregs_26__18_,
         decode_regfile_intregs_26__19_, decode_regfile_intregs_26__20_,
         decode_regfile_intregs_26__21_, decode_regfile_intregs_26__22_,
         decode_regfile_intregs_26__23_, decode_regfile_intregs_26__24_,
         decode_regfile_intregs_26__25_, decode_regfile_intregs_26__26_,
         decode_regfile_intregs_26__27_, decode_regfile_intregs_26__28_,
         decode_regfile_intregs_26__29_, decode_regfile_intregs_26__30_,
         decode_regfile_intregs_26__31_, decode_regfile_intregs_27__0_,
         decode_regfile_intregs_27__1_, decode_regfile_intregs_27__2_,
         decode_regfile_intregs_27__3_, decode_regfile_intregs_27__4_,
         decode_regfile_intregs_27__5_, decode_regfile_intregs_27__6_,
         decode_regfile_intregs_27__7_, decode_regfile_intregs_27__8_,
         decode_regfile_intregs_27__9_, decode_regfile_intregs_27__10_,
         decode_regfile_intregs_27__11_, decode_regfile_intregs_27__12_,
         decode_regfile_intregs_27__13_, decode_regfile_intregs_27__14_,
         decode_regfile_intregs_27__15_, decode_regfile_intregs_27__16_,
         decode_regfile_intregs_27__17_, decode_regfile_intregs_27__18_,
         decode_regfile_intregs_27__19_, decode_regfile_intregs_27__20_,
         decode_regfile_intregs_27__21_, decode_regfile_intregs_27__22_,
         decode_regfile_intregs_27__23_, decode_regfile_intregs_27__24_,
         decode_regfile_intregs_27__25_, decode_regfile_intregs_27__26_,
         decode_regfile_intregs_27__27_, decode_regfile_intregs_27__28_,
         decode_regfile_intregs_27__29_, decode_regfile_intregs_27__30_,
         decode_regfile_intregs_27__31_, decode_regfile_intregs_28__0_,
         decode_regfile_intregs_28__1_, decode_regfile_intregs_28__2_,
         decode_regfile_intregs_28__3_, decode_regfile_intregs_28__4_,
         decode_regfile_intregs_28__5_, decode_regfile_intregs_28__6_,
         decode_regfile_intregs_28__7_, decode_regfile_intregs_28__8_,
         decode_regfile_intregs_28__9_, decode_regfile_intregs_28__10_,
         decode_regfile_intregs_28__11_, decode_regfile_intregs_28__12_,
         decode_regfile_intregs_28__13_, decode_regfile_intregs_28__14_,
         decode_regfile_intregs_28__15_, decode_regfile_intregs_28__16_,
         decode_regfile_intregs_28__17_, decode_regfile_intregs_28__18_,
         decode_regfile_intregs_28__19_, decode_regfile_intregs_28__20_,
         decode_regfile_intregs_28__21_, decode_regfile_intregs_28__22_,
         decode_regfile_intregs_28__23_, decode_regfile_intregs_28__24_,
         decode_regfile_intregs_28__25_, decode_regfile_intregs_28__26_,
         decode_regfile_intregs_28__27_, decode_regfile_intregs_28__28_,
         decode_regfile_intregs_28__29_, decode_regfile_intregs_28__30_,
         decode_regfile_intregs_28__31_, decode_regfile_intregs_29__0_,
         decode_regfile_intregs_29__1_, decode_regfile_intregs_29__2_,
         decode_regfile_intregs_29__3_, decode_regfile_intregs_29__4_,
         decode_regfile_intregs_29__5_, decode_regfile_intregs_29__6_,
         decode_regfile_intregs_29__7_, decode_regfile_intregs_29__8_,
         decode_regfile_intregs_29__9_, decode_regfile_intregs_29__10_,
         decode_regfile_intregs_29__11_, decode_regfile_intregs_29__12_,
         decode_regfile_intregs_29__13_, decode_regfile_intregs_29__14_,
         decode_regfile_intregs_29__15_, decode_regfile_intregs_29__16_,
         decode_regfile_intregs_29__17_, decode_regfile_intregs_29__18_,
         decode_regfile_intregs_29__19_, decode_regfile_intregs_29__20_,
         decode_regfile_intregs_29__21_, decode_regfile_intregs_29__22_,
         decode_regfile_intregs_29__23_, decode_regfile_intregs_29__24_,
         decode_regfile_intregs_29__25_, decode_regfile_intregs_29__26_,
         decode_regfile_intregs_29__27_, decode_regfile_intregs_29__28_,
         decode_regfile_intregs_29__29_, decode_regfile_intregs_29__30_,
         decode_regfile_intregs_29__31_, decode_regfile_intregs_30__0_,
         decode_regfile_intregs_30__1_, decode_regfile_intregs_30__2_,
         decode_regfile_intregs_30__3_, decode_regfile_intregs_30__4_,
         decode_regfile_intregs_30__5_, decode_regfile_intregs_30__6_,
         decode_regfile_intregs_30__7_, decode_regfile_intregs_30__8_,
         decode_regfile_intregs_30__9_, decode_regfile_intregs_30__10_,
         decode_regfile_intregs_30__11_, decode_regfile_intregs_30__12_,
         decode_regfile_intregs_30__13_, decode_regfile_intregs_30__14_,
         decode_regfile_intregs_30__15_, decode_regfile_intregs_30__16_,
         decode_regfile_intregs_30__17_, decode_regfile_intregs_30__18_,
         decode_regfile_intregs_30__19_, decode_regfile_intregs_30__20_,
         decode_regfile_intregs_30__21_, decode_regfile_intregs_30__22_,
         decode_regfile_intregs_30__23_, decode_regfile_intregs_30__24_,
         decode_regfile_intregs_30__25_, decode_regfile_intregs_30__26_,
         decode_regfile_intregs_30__27_, decode_regfile_intregs_30__28_,
         decode_regfile_intregs_30__29_, decode_regfile_intregs_30__30_,
         decode_regfile_intregs_30__31_, decode_regfile_intregs_31__0_,
         decode_regfile_intregs_31__1_, decode_regfile_intregs_31__2_,
         decode_regfile_intregs_31__3_, decode_regfile_intregs_31__4_,
         decode_regfile_intregs_31__5_, decode_regfile_intregs_31__6_,
         decode_regfile_intregs_31__7_, decode_regfile_intregs_31__8_,
         decode_regfile_intregs_31__9_, decode_regfile_intregs_31__10_,
         decode_regfile_intregs_31__11_, decode_regfile_intregs_31__12_,
         decode_regfile_intregs_31__13_, decode_regfile_intregs_31__14_,
         decode_regfile_intregs_31__15_, decode_regfile_intregs_31__16_,
         decode_regfile_intregs_31__17_, decode_regfile_intregs_31__18_,
         decode_regfile_intregs_31__19_, decode_regfile_intregs_31__20_,
         decode_regfile_intregs_31__21_, decode_regfile_intregs_31__22_,
         decode_regfile_intregs_31__23_, decode_regfile_intregs_31__24_,
         decode_regfile_intregs_31__25_, decode_regfile_intregs_31__26_,
         decode_regfile_intregs_31__27_, decode_regfile_intregs_31__28_,
         decode_regfile_intregs_31__29_, decode_regfile_intregs_31__30_,
         decode_regfile_intregs_31__31_, decode_regfile_fpregs_0__0_,
         decode_regfile_fpregs_0__1_, decode_regfile_fpregs_0__2_,
         decode_regfile_fpregs_0__3_, decode_regfile_fpregs_0__4_,
         decode_regfile_fpregs_0__5_, decode_regfile_fpregs_0__6_,
         decode_regfile_fpregs_0__7_, decode_regfile_fpregs_0__8_,
         decode_regfile_fpregs_0__9_, decode_regfile_fpregs_0__10_,
         decode_regfile_fpregs_0__11_, decode_regfile_fpregs_0__12_,
         decode_regfile_fpregs_0__13_, decode_regfile_fpregs_0__14_,
         decode_regfile_fpregs_0__15_, decode_regfile_fpregs_0__16_,
         decode_regfile_fpregs_0__17_, decode_regfile_fpregs_0__18_,
         decode_regfile_fpregs_0__19_, decode_regfile_fpregs_0__20_,
         decode_regfile_fpregs_0__21_, decode_regfile_fpregs_0__22_,
         decode_regfile_fpregs_0__23_, decode_regfile_fpregs_0__24_,
         decode_regfile_fpregs_0__25_, decode_regfile_fpregs_0__26_,
         decode_regfile_fpregs_0__27_, decode_regfile_fpregs_0__28_,
         decode_regfile_fpregs_0__29_, decode_regfile_fpregs_0__30_,
         decode_regfile_fpregs_0__31_, decode_regfile_fpregs_1__0_,
         decode_regfile_fpregs_1__1_, decode_regfile_fpregs_1__2_,
         decode_regfile_fpregs_1__3_, decode_regfile_fpregs_1__4_,
         decode_regfile_fpregs_1__5_, decode_regfile_fpregs_1__6_,
         decode_regfile_fpregs_1__7_, decode_regfile_fpregs_1__8_,
         decode_regfile_fpregs_1__9_, decode_regfile_fpregs_1__10_,
         decode_regfile_fpregs_1__11_, decode_regfile_fpregs_1__12_,
         decode_regfile_fpregs_1__13_, decode_regfile_fpregs_1__14_,
         decode_regfile_fpregs_1__15_, decode_regfile_fpregs_1__16_,
         decode_regfile_fpregs_1__17_, decode_regfile_fpregs_1__18_,
         decode_regfile_fpregs_1__19_, decode_regfile_fpregs_1__20_,
         decode_regfile_fpregs_1__21_, decode_regfile_fpregs_1__22_,
         decode_regfile_fpregs_1__23_, decode_regfile_fpregs_1__24_,
         decode_regfile_fpregs_1__25_, decode_regfile_fpregs_1__26_,
         decode_regfile_fpregs_1__27_, decode_regfile_fpregs_1__28_,
         decode_regfile_fpregs_1__29_, decode_regfile_fpregs_1__30_,
         decode_regfile_fpregs_1__31_, decode_regfile_fpregs_2__0_,
         decode_regfile_fpregs_2__1_, decode_regfile_fpregs_2__2_,
         decode_regfile_fpregs_2__3_, decode_regfile_fpregs_2__4_,
         decode_regfile_fpregs_2__5_, decode_regfile_fpregs_2__6_,
         decode_regfile_fpregs_2__7_, decode_regfile_fpregs_2__8_,
         decode_regfile_fpregs_2__9_, decode_regfile_fpregs_2__10_,
         decode_regfile_fpregs_2__11_, decode_regfile_fpregs_2__12_,
         decode_regfile_fpregs_2__13_, decode_regfile_fpregs_2__14_,
         decode_regfile_fpregs_2__15_, decode_regfile_fpregs_2__16_,
         decode_regfile_fpregs_2__17_, decode_regfile_fpregs_2__18_,
         decode_regfile_fpregs_2__19_, decode_regfile_fpregs_2__20_,
         decode_regfile_fpregs_2__21_, decode_regfile_fpregs_2__22_,
         decode_regfile_fpregs_2__23_, decode_regfile_fpregs_2__24_,
         decode_regfile_fpregs_2__25_, decode_regfile_fpregs_2__26_,
         decode_regfile_fpregs_2__27_, decode_regfile_fpregs_2__28_,
         decode_regfile_fpregs_2__29_, decode_regfile_fpregs_2__30_,
         decode_regfile_fpregs_2__31_, decode_regfile_fpregs_3__0_,
         decode_regfile_fpregs_3__1_, decode_regfile_fpregs_3__2_,
         decode_regfile_fpregs_3__3_, decode_regfile_fpregs_3__4_,
         decode_regfile_fpregs_3__5_, decode_regfile_fpregs_3__6_,
         decode_regfile_fpregs_3__7_, decode_regfile_fpregs_3__8_,
         decode_regfile_fpregs_3__9_, decode_regfile_fpregs_3__10_,
         decode_regfile_fpregs_3__11_, decode_regfile_fpregs_3__12_,
         decode_regfile_fpregs_3__13_, decode_regfile_fpregs_3__14_,
         decode_regfile_fpregs_3__15_, decode_regfile_fpregs_3__16_,
         decode_regfile_fpregs_3__17_, decode_regfile_fpregs_3__18_,
         decode_regfile_fpregs_3__19_, decode_regfile_fpregs_3__20_,
         decode_regfile_fpregs_3__21_, decode_regfile_fpregs_3__22_,
         decode_regfile_fpregs_3__23_, decode_regfile_fpregs_3__24_,
         decode_regfile_fpregs_3__25_, decode_regfile_fpregs_3__26_,
         decode_regfile_fpregs_3__27_, decode_regfile_fpregs_3__28_,
         decode_regfile_fpregs_3__29_, decode_regfile_fpregs_3__30_,
         decode_regfile_fpregs_3__31_, decode_regfile_fpregs_4__0_,
         decode_regfile_fpregs_4__1_, decode_regfile_fpregs_4__2_,
         decode_regfile_fpregs_4__3_, decode_regfile_fpregs_4__4_,
         decode_regfile_fpregs_4__5_, decode_regfile_fpregs_4__6_,
         decode_regfile_fpregs_4__7_, decode_regfile_fpregs_4__8_,
         decode_regfile_fpregs_4__9_, decode_regfile_fpregs_4__10_,
         decode_regfile_fpregs_4__11_, decode_regfile_fpregs_4__12_,
         decode_regfile_fpregs_4__13_, decode_regfile_fpregs_4__14_,
         decode_regfile_fpregs_4__15_, decode_regfile_fpregs_4__16_,
         decode_regfile_fpregs_4__17_, decode_regfile_fpregs_4__18_,
         decode_regfile_fpregs_4__19_, decode_regfile_fpregs_4__20_,
         decode_regfile_fpregs_4__21_, decode_regfile_fpregs_4__22_,
         decode_regfile_fpregs_4__23_, decode_regfile_fpregs_4__24_,
         decode_regfile_fpregs_4__25_, decode_regfile_fpregs_4__26_,
         decode_regfile_fpregs_4__27_, decode_regfile_fpregs_4__28_,
         decode_regfile_fpregs_4__29_, decode_regfile_fpregs_4__30_,
         decode_regfile_fpregs_4__31_, decode_regfile_fpregs_5__0_,
         decode_regfile_fpregs_5__1_, decode_regfile_fpregs_5__2_,
         decode_regfile_fpregs_5__3_, decode_regfile_fpregs_5__4_,
         decode_regfile_fpregs_5__5_, decode_regfile_fpregs_5__6_,
         decode_regfile_fpregs_5__7_, decode_regfile_fpregs_5__8_,
         decode_regfile_fpregs_5__9_, decode_regfile_fpregs_5__10_,
         decode_regfile_fpregs_5__11_, decode_regfile_fpregs_5__12_,
         decode_regfile_fpregs_5__13_, decode_regfile_fpregs_5__14_,
         decode_regfile_fpregs_5__15_, decode_regfile_fpregs_5__16_,
         decode_regfile_fpregs_5__17_, decode_regfile_fpregs_5__18_,
         decode_regfile_fpregs_5__19_, decode_regfile_fpregs_5__20_,
         decode_regfile_fpregs_5__21_, decode_regfile_fpregs_5__22_,
         decode_regfile_fpregs_5__23_, decode_regfile_fpregs_5__24_,
         decode_regfile_fpregs_5__25_, decode_regfile_fpregs_5__26_,
         decode_regfile_fpregs_5__27_, decode_regfile_fpregs_5__28_,
         decode_regfile_fpregs_5__29_, decode_regfile_fpregs_5__30_,
         decode_regfile_fpregs_5__31_, decode_regfile_fpregs_6__0_,
         decode_regfile_fpregs_6__1_, decode_regfile_fpregs_6__2_,
         decode_regfile_fpregs_6__3_, decode_regfile_fpregs_6__4_,
         decode_regfile_fpregs_6__5_, decode_regfile_fpregs_6__6_,
         decode_regfile_fpregs_6__7_, decode_regfile_fpregs_6__8_,
         decode_regfile_fpregs_6__9_, decode_regfile_fpregs_6__10_,
         decode_regfile_fpregs_6__11_, decode_regfile_fpregs_6__12_,
         decode_regfile_fpregs_6__13_, decode_regfile_fpregs_6__14_,
         decode_regfile_fpregs_6__15_, decode_regfile_fpregs_6__16_,
         decode_regfile_fpregs_6__17_, decode_regfile_fpregs_6__18_,
         decode_regfile_fpregs_6__19_, decode_regfile_fpregs_6__20_,
         decode_regfile_fpregs_6__21_, decode_regfile_fpregs_6__22_,
         decode_regfile_fpregs_6__23_, decode_regfile_fpregs_6__24_,
         decode_regfile_fpregs_6__25_, decode_regfile_fpregs_6__26_,
         decode_regfile_fpregs_6__27_, decode_regfile_fpregs_6__28_,
         decode_regfile_fpregs_6__29_, decode_regfile_fpregs_6__30_,
         decode_regfile_fpregs_6__31_, decode_regfile_fpregs_7__0_,
         decode_regfile_fpregs_7__1_, decode_regfile_fpregs_7__2_,
         decode_regfile_fpregs_7__3_, decode_regfile_fpregs_7__4_,
         decode_regfile_fpregs_7__5_, decode_regfile_fpregs_7__6_,
         decode_regfile_fpregs_7__7_, decode_regfile_fpregs_7__8_,
         decode_regfile_fpregs_7__9_, decode_regfile_fpregs_7__10_,
         decode_regfile_fpregs_7__11_, decode_regfile_fpregs_7__12_,
         decode_regfile_fpregs_7__13_, decode_regfile_fpregs_7__14_,
         decode_regfile_fpregs_7__15_, decode_regfile_fpregs_7__16_,
         decode_regfile_fpregs_7__17_, decode_regfile_fpregs_7__18_,
         decode_regfile_fpregs_7__19_, decode_regfile_fpregs_7__20_,
         decode_regfile_fpregs_7__21_, decode_regfile_fpregs_7__22_,
         decode_regfile_fpregs_7__23_, decode_regfile_fpregs_7__24_,
         decode_regfile_fpregs_7__25_, decode_regfile_fpregs_7__26_,
         decode_regfile_fpregs_7__27_, decode_regfile_fpregs_7__28_,
         decode_regfile_fpregs_7__29_, decode_regfile_fpregs_7__30_,
         decode_regfile_fpregs_7__31_, decode_regfile_fpregs_8__0_,
         decode_regfile_fpregs_8__1_, decode_regfile_fpregs_8__2_,
         decode_regfile_fpregs_8__3_, decode_regfile_fpregs_8__4_,
         decode_regfile_fpregs_8__5_, decode_regfile_fpregs_8__6_,
         decode_regfile_fpregs_8__7_, decode_regfile_fpregs_8__8_,
         decode_regfile_fpregs_8__9_, decode_regfile_fpregs_8__10_,
         decode_regfile_fpregs_8__11_, decode_regfile_fpregs_8__12_,
         decode_regfile_fpregs_8__13_, decode_regfile_fpregs_8__14_,
         decode_regfile_fpregs_8__15_, decode_regfile_fpregs_8__16_,
         decode_regfile_fpregs_8__17_, decode_regfile_fpregs_8__18_,
         decode_regfile_fpregs_8__19_, decode_regfile_fpregs_8__20_,
         decode_regfile_fpregs_8__21_, decode_regfile_fpregs_8__22_,
         decode_regfile_fpregs_8__23_, decode_regfile_fpregs_8__24_,
         decode_regfile_fpregs_8__25_, decode_regfile_fpregs_8__26_,
         decode_regfile_fpregs_8__27_, decode_regfile_fpregs_8__28_,
         decode_regfile_fpregs_8__29_, decode_regfile_fpregs_8__30_,
         decode_regfile_fpregs_8__31_, decode_regfile_fpregs_9__0_,
         decode_regfile_fpregs_9__1_, decode_regfile_fpregs_9__2_,
         decode_regfile_fpregs_9__3_, decode_regfile_fpregs_9__4_,
         decode_regfile_fpregs_9__5_, decode_regfile_fpregs_9__6_,
         decode_regfile_fpregs_9__7_, decode_regfile_fpregs_9__8_,
         decode_regfile_fpregs_9__9_, decode_regfile_fpregs_9__10_,
         decode_regfile_fpregs_9__11_, decode_regfile_fpregs_9__12_,
         decode_regfile_fpregs_9__13_, decode_regfile_fpregs_9__14_,
         decode_regfile_fpregs_9__15_, decode_regfile_fpregs_9__16_,
         decode_regfile_fpregs_9__17_, decode_regfile_fpregs_9__18_,
         decode_regfile_fpregs_9__19_, decode_regfile_fpregs_9__20_,
         decode_regfile_fpregs_9__21_, decode_regfile_fpregs_9__22_,
         decode_regfile_fpregs_9__23_, decode_regfile_fpregs_9__24_,
         decode_regfile_fpregs_9__25_, decode_regfile_fpregs_9__26_,
         decode_regfile_fpregs_9__27_, decode_regfile_fpregs_9__28_,
         decode_regfile_fpregs_9__29_, decode_regfile_fpregs_9__30_,
         decode_regfile_fpregs_9__31_, decode_regfile_fpregs_10__0_,
         decode_regfile_fpregs_10__1_, decode_regfile_fpregs_10__2_,
         decode_regfile_fpregs_10__3_, decode_regfile_fpregs_10__4_,
         decode_regfile_fpregs_10__5_, decode_regfile_fpregs_10__6_,
         decode_regfile_fpregs_10__7_, decode_regfile_fpregs_10__8_,
         decode_regfile_fpregs_10__9_, decode_regfile_fpregs_10__10_,
         decode_regfile_fpregs_10__11_, decode_regfile_fpregs_10__12_,
         decode_regfile_fpregs_10__13_, decode_regfile_fpregs_10__14_,
         decode_regfile_fpregs_10__15_, decode_regfile_fpregs_10__16_,
         decode_regfile_fpregs_10__17_, decode_regfile_fpregs_10__18_,
         decode_regfile_fpregs_10__19_, decode_regfile_fpregs_10__20_,
         decode_regfile_fpregs_10__21_, decode_regfile_fpregs_10__22_,
         decode_regfile_fpregs_10__23_, decode_regfile_fpregs_10__24_,
         decode_regfile_fpregs_10__25_, decode_regfile_fpregs_10__26_,
         decode_regfile_fpregs_10__27_, decode_regfile_fpregs_10__28_,
         decode_regfile_fpregs_10__29_, decode_regfile_fpregs_10__30_,
         decode_regfile_fpregs_10__31_, decode_regfile_fpregs_11__0_,
         decode_regfile_fpregs_11__1_, decode_regfile_fpregs_11__2_,
         decode_regfile_fpregs_11__3_, decode_regfile_fpregs_11__4_,
         decode_regfile_fpregs_11__5_, decode_regfile_fpregs_11__6_,
         decode_regfile_fpregs_11__7_, decode_regfile_fpregs_11__8_,
         decode_regfile_fpregs_11__9_, decode_regfile_fpregs_11__10_,
         decode_regfile_fpregs_11__11_, decode_regfile_fpregs_11__12_,
         decode_regfile_fpregs_11__13_, decode_regfile_fpregs_11__14_,
         decode_regfile_fpregs_11__15_, decode_regfile_fpregs_11__16_,
         decode_regfile_fpregs_11__17_, decode_regfile_fpregs_11__18_,
         decode_regfile_fpregs_11__19_, decode_regfile_fpregs_11__20_,
         decode_regfile_fpregs_11__21_, decode_regfile_fpregs_11__22_,
         decode_regfile_fpregs_11__23_, decode_regfile_fpregs_11__24_,
         decode_regfile_fpregs_11__25_, decode_regfile_fpregs_11__26_,
         decode_regfile_fpregs_11__27_, decode_regfile_fpregs_11__28_,
         decode_regfile_fpregs_11__29_, decode_regfile_fpregs_11__30_,
         decode_regfile_fpregs_11__31_, decode_regfile_fpregs_12__0_,
         decode_regfile_fpregs_12__1_, decode_regfile_fpregs_12__2_,
         decode_regfile_fpregs_12__3_, decode_regfile_fpregs_12__4_,
         decode_regfile_fpregs_12__5_, decode_regfile_fpregs_12__6_,
         decode_regfile_fpregs_12__7_, decode_regfile_fpregs_12__8_,
         decode_regfile_fpregs_12__9_, decode_regfile_fpregs_12__10_,
         decode_regfile_fpregs_12__11_, decode_regfile_fpregs_12__12_,
         decode_regfile_fpregs_12__13_, decode_regfile_fpregs_12__14_,
         decode_regfile_fpregs_12__15_, decode_regfile_fpregs_12__16_,
         decode_regfile_fpregs_12__17_, decode_regfile_fpregs_12__18_,
         decode_regfile_fpregs_12__19_, decode_regfile_fpregs_12__20_,
         decode_regfile_fpregs_12__21_, decode_regfile_fpregs_12__22_,
         decode_regfile_fpregs_12__23_, decode_regfile_fpregs_12__24_,
         decode_regfile_fpregs_12__25_, decode_regfile_fpregs_12__26_,
         decode_regfile_fpregs_12__27_, decode_regfile_fpregs_12__28_,
         decode_regfile_fpregs_12__29_, decode_regfile_fpregs_12__30_,
         decode_regfile_fpregs_12__31_, decode_regfile_fpregs_13__0_,
         decode_regfile_fpregs_13__1_, decode_regfile_fpregs_13__2_,
         decode_regfile_fpregs_13__3_, decode_regfile_fpregs_13__4_,
         decode_regfile_fpregs_13__5_, decode_regfile_fpregs_13__6_,
         decode_regfile_fpregs_13__7_, decode_regfile_fpregs_13__8_,
         decode_regfile_fpregs_13__9_, decode_regfile_fpregs_13__10_,
         decode_regfile_fpregs_13__11_, decode_regfile_fpregs_13__12_,
         decode_regfile_fpregs_13__13_, decode_regfile_fpregs_13__14_,
         decode_regfile_fpregs_13__15_, decode_regfile_fpregs_13__16_,
         decode_regfile_fpregs_13__17_, decode_regfile_fpregs_13__18_,
         decode_regfile_fpregs_13__19_, decode_regfile_fpregs_13__20_,
         decode_regfile_fpregs_13__21_, decode_regfile_fpregs_13__22_,
         decode_regfile_fpregs_13__23_, decode_regfile_fpregs_13__24_,
         decode_regfile_fpregs_13__25_, decode_regfile_fpregs_13__26_,
         decode_regfile_fpregs_13__27_, decode_regfile_fpregs_13__28_,
         decode_regfile_fpregs_13__29_, decode_regfile_fpregs_13__30_,
         decode_regfile_fpregs_13__31_, decode_regfile_fpregs_14__0_,
         decode_regfile_fpregs_14__1_, decode_regfile_fpregs_14__2_,
         decode_regfile_fpregs_14__3_, decode_regfile_fpregs_14__4_,
         decode_regfile_fpregs_14__5_, decode_regfile_fpregs_14__6_,
         decode_regfile_fpregs_14__7_, decode_regfile_fpregs_14__8_,
         decode_regfile_fpregs_14__9_, decode_regfile_fpregs_14__10_,
         decode_regfile_fpregs_14__11_, decode_regfile_fpregs_14__12_,
         decode_regfile_fpregs_14__13_, decode_regfile_fpregs_14__14_,
         decode_regfile_fpregs_14__15_, decode_regfile_fpregs_14__16_,
         decode_regfile_fpregs_14__17_, decode_regfile_fpregs_14__18_,
         decode_regfile_fpregs_14__19_, decode_regfile_fpregs_14__20_,
         decode_regfile_fpregs_14__21_, decode_regfile_fpregs_14__22_,
         decode_regfile_fpregs_14__23_, decode_regfile_fpregs_14__24_,
         decode_regfile_fpregs_14__25_, decode_regfile_fpregs_14__26_,
         decode_regfile_fpregs_14__27_, decode_regfile_fpregs_14__28_,
         decode_regfile_fpregs_14__29_, decode_regfile_fpregs_14__30_,
         decode_regfile_fpregs_14__31_, decode_regfile_fpregs_15__0_,
         decode_regfile_fpregs_15__1_, decode_regfile_fpregs_15__2_,
         decode_regfile_fpregs_15__3_, decode_regfile_fpregs_15__4_,
         decode_regfile_fpregs_15__5_, decode_regfile_fpregs_15__6_,
         decode_regfile_fpregs_15__7_, decode_regfile_fpregs_15__8_,
         decode_regfile_fpregs_15__9_, decode_regfile_fpregs_15__10_,
         decode_regfile_fpregs_15__11_, decode_regfile_fpregs_15__12_,
         decode_regfile_fpregs_15__13_, decode_regfile_fpregs_15__14_,
         decode_regfile_fpregs_15__15_, decode_regfile_fpregs_15__16_,
         decode_regfile_fpregs_15__17_, decode_regfile_fpregs_15__18_,
         decode_regfile_fpregs_15__19_, decode_regfile_fpregs_15__20_,
         decode_regfile_fpregs_15__21_, decode_regfile_fpregs_15__22_,
         decode_regfile_fpregs_15__23_, decode_regfile_fpregs_15__24_,
         decode_regfile_fpregs_15__25_, decode_regfile_fpregs_15__26_,
         decode_regfile_fpregs_15__27_, decode_regfile_fpregs_15__28_,
         decode_regfile_fpregs_15__29_, decode_regfile_fpregs_15__30_,
         decode_regfile_fpregs_15__31_, decode_regfile_fpregs_16__0_,
         decode_regfile_fpregs_16__1_, decode_regfile_fpregs_16__2_,
         decode_regfile_fpregs_16__3_, decode_regfile_fpregs_16__4_,
         decode_regfile_fpregs_16__5_, decode_regfile_fpregs_16__6_,
         decode_regfile_fpregs_16__7_, decode_regfile_fpregs_16__8_,
         decode_regfile_fpregs_16__9_, decode_regfile_fpregs_16__10_,
         decode_regfile_fpregs_16__11_, decode_regfile_fpregs_16__12_,
         decode_regfile_fpregs_16__13_, decode_regfile_fpregs_16__14_,
         decode_regfile_fpregs_16__15_, decode_regfile_fpregs_16__16_,
         decode_regfile_fpregs_16__17_, decode_regfile_fpregs_16__18_,
         decode_regfile_fpregs_16__19_, decode_regfile_fpregs_16__20_,
         decode_regfile_fpregs_16__21_, decode_regfile_fpregs_16__22_,
         decode_regfile_fpregs_16__23_, decode_regfile_fpregs_16__24_,
         decode_regfile_fpregs_16__25_, decode_regfile_fpregs_16__26_,
         decode_regfile_fpregs_16__27_, decode_regfile_fpregs_16__28_,
         decode_regfile_fpregs_16__29_, decode_regfile_fpregs_16__30_,
         decode_regfile_fpregs_16__31_, decode_regfile_fpregs_17__0_,
         decode_regfile_fpregs_17__1_, decode_regfile_fpregs_17__2_,
         decode_regfile_fpregs_17__3_, decode_regfile_fpregs_17__4_,
         decode_regfile_fpregs_17__5_, decode_regfile_fpregs_17__6_,
         decode_regfile_fpregs_17__7_, decode_regfile_fpregs_17__8_,
         decode_regfile_fpregs_17__9_, decode_regfile_fpregs_17__10_,
         decode_regfile_fpregs_17__11_, decode_regfile_fpregs_17__12_,
         decode_regfile_fpregs_17__13_, decode_regfile_fpregs_17__14_,
         decode_regfile_fpregs_17__15_, decode_regfile_fpregs_17__16_,
         decode_regfile_fpregs_17__17_, decode_regfile_fpregs_17__18_,
         decode_regfile_fpregs_17__19_, decode_regfile_fpregs_17__20_,
         decode_regfile_fpregs_17__21_, decode_regfile_fpregs_17__22_,
         decode_regfile_fpregs_17__23_, decode_regfile_fpregs_17__24_,
         decode_regfile_fpregs_17__25_, decode_regfile_fpregs_17__26_,
         decode_regfile_fpregs_17__27_, decode_regfile_fpregs_17__28_,
         decode_regfile_fpregs_17__29_, decode_regfile_fpregs_17__30_,
         decode_regfile_fpregs_17__31_, decode_regfile_fpregs_18__0_,
         decode_regfile_fpregs_18__1_, decode_regfile_fpregs_18__2_,
         decode_regfile_fpregs_18__3_, decode_regfile_fpregs_18__4_,
         decode_regfile_fpregs_18__5_, decode_regfile_fpregs_18__6_,
         decode_regfile_fpregs_18__7_, decode_regfile_fpregs_18__8_,
         decode_regfile_fpregs_18__9_, decode_regfile_fpregs_18__10_,
         decode_regfile_fpregs_18__11_, decode_regfile_fpregs_18__12_,
         decode_regfile_fpregs_18__13_, decode_regfile_fpregs_18__14_,
         decode_regfile_fpregs_18__15_, decode_regfile_fpregs_18__16_,
         decode_regfile_fpregs_18__17_, decode_regfile_fpregs_18__18_,
         decode_regfile_fpregs_18__19_, decode_regfile_fpregs_18__20_,
         decode_regfile_fpregs_18__21_, decode_regfile_fpregs_18__22_,
         decode_regfile_fpregs_18__23_, decode_regfile_fpregs_18__24_,
         decode_regfile_fpregs_18__25_, decode_regfile_fpregs_18__26_,
         decode_regfile_fpregs_18__27_, decode_regfile_fpregs_18__28_,
         decode_regfile_fpregs_18__29_, decode_regfile_fpregs_18__30_,
         decode_regfile_fpregs_18__31_, decode_regfile_fpregs_19__0_,
         decode_regfile_fpregs_19__1_, decode_regfile_fpregs_19__2_,
         decode_regfile_fpregs_19__3_, decode_regfile_fpregs_19__4_,
         decode_regfile_fpregs_19__5_, decode_regfile_fpregs_19__6_,
         decode_regfile_fpregs_19__7_, decode_regfile_fpregs_19__8_,
         decode_regfile_fpregs_19__9_, decode_regfile_fpregs_19__10_,
         decode_regfile_fpregs_19__11_, decode_regfile_fpregs_19__12_,
         decode_regfile_fpregs_19__13_, decode_regfile_fpregs_19__14_,
         decode_regfile_fpregs_19__15_, decode_regfile_fpregs_19__16_,
         decode_regfile_fpregs_19__17_, decode_regfile_fpregs_19__18_,
         decode_regfile_fpregs_19__19_, decode_regfile_fpregs_19__20_,
         decode_regfile_fpregs_19__21_, decode_regfile_fpregs_19__22_,
         decode_regfile_fpregs_19__23_, decode_regfile_fpregs_19__24_,
         decode_regfile_fpregs_19__25_, decode_regfile_fpregs_19__26_,
         decode_regfile_fpregs_19__27_, decode_regfile_fpregs_19__28_,
         decode_regfile_fpregs_19__29_, decode_regfile_fpregs_19__30_,
         decode_regfile_fpregs_19__31_, decode_regfile_fpregs_20__0_,
         decode_regfile_fpregs_20__1_, decode_regfile_fpregs_20__2_,
         decode_regfile_fpregs_20__3_, decode_regfile_fpregs_20__4_,
         decode_regfile_fpregs_20__5_, decode_regfile_fpregs_20__6_,
         decode_regfile_fpregs_20__7_, decode_regfile_fpregs_20__8_,
         decode_regfile_fpregs_20__9_, decode_regfile_fpregs_20__10_,
         decode_regfile_fpregs_20__11_, decode_regfile_fpregs_20__12_,
         decode_regfile_fpregs_20__13_, decode_regfile_fpregs_20__14_,
         decode_regfile_fpregs_20__15_, decode_regfile_fpregs_20__16_,
         decode_regfile_fpregs_20__17_, decode_regfile_fpregs_20__18_,
         decode_regfile_fpregs_20__19_, decode_regfile_fpregs_20__20_,
         decode_regfile_fpregs_20__21_, decode_regfile_fpregs_20__22_,
         decode_regfile_fpregs_20__23_, decode_regfile_fpregs_20__24_,
         decode_regfile_fpregs_20__25_, decode_regfile_fpregs_20__26_,
         decode_regfile_fpregs_20__27_, decode_regfile_fpregs_20__28_,
         decode_regfile_fpregs_20__29_, decode_regfile_fpregs_20__30_,
         decode_regfile_fpregs_20__31_, decode_regfile_fpregs_21__0_,
         decode_regfile_fpregs_21__1_, decode_regfile_fpregs_21__2_,
         decode_regfile_fpregs_21__3_, decode_regfile_fpregs_21__4_,
         decode_regfile_fpregs_21__5_, decode_regfile_fpregs_21__6_,
         decode_regfile_fpregs_21__7_, decode_regfile_fpregs_21__8_,
         decode_regfile_fpregs_21__9_, decode_regfile_fpregs_21__10_,
         decode_regfile_fpregs_21__11_, decode_regfile_fpregs_21__12_,
         decode_regfile_fpregs_21__13_, decode_regfile_fpregs_21__14_,
         decode_regfile_fpregs_21__15_, decode_regfile_fpregs_21__16_,
         decode_regfile_fpregs_21__17_, decode_regfile_fpregs_21__18_,
         decode_regfile_fpregs_21__19_, decode_regfile_fpregs_21__20_,
         decode_regfile_fpregs_21__21_, decode_regfile_fpregs_21__22_,
         decode_regfile_fpregs_21__23_, decode_regfile_fpregs_21__24_,
         decode_regfile_fpregs_21__25_, decode_regfile_fpregs_21__26_,
         decode_regfile_fpregs_21__27_, decode_regfile_fpregs_21__28_,
         decode_regfile_fpregs_21__29_, decode_regfile_fpregs_21__30_,
         decode_regfile_fpregs_21__31_, decode_regfile_fpregs_22__0_,
         decode_regfile_fpregs_22__1_, decode_regfile_fpregs_22__2_,
         decode_regfile_fpregs_22__3_, decode_regfile_fpregs_22__4_,
         decode_regfile_fpregs_22__5_, decode_regfile_fpregs_22__6_,
         decode_regfile_fpregs_22__7_, decode_regfile_fpregs_22__8_,
         decode_regfile_fpregs_22__9_, decode_regfile_fpregs_22__10_,
         decode_regfile_fpregs_22__11_, decode_regfile_fpregs_22__12_,
         decode_regfile_fpregs_22__13_, decode_regfile_fpregs_22__14_,
         decode_regfile_fpregs_22__15_, decode_regfile_fpregs_22__16_,
         decode_regfile_fpregs_22__17_, decode_regfile_fpregs_22__18_,
         decode_regfile_fpregs_22__19_, decode_regfile_fpregs_22__20_,
         decode_regfile_fpregs_22__21_, decode_regfile_fpregs_22__22_,
         decode_regfile_fpregs_22__23_, decode_regfile_fpregs_22__24_,
         decode_regfile_fpregs_22__25_, decode_regfile_fpregs_22__26_,
         decode_regfile_fpregs_22__27_, decode_regfile_fpregs_22__28_,
         decode_regfile_fpregs_22__29_, decode_regfile_fpregs_22__30_,
         decode_regfile_fpregs_22__31_, decode_regfile_fpregs_23__0_,
         decode_regfile_fpregs_23__1_, decode_regfile_fpregs_23__2_,
         decode_regfile_fpregs_23__3_, decode_regfile_fpregs_23__4_,
         decode_regfile_fpregs_23__5_, decode_regfile_fpregs_23__6_,
         decode_regfile_fpregs_23__7_, decode_regfile_fpregs_23__8_,
         decode_regfile_fpregs_23__9_, decode_regfile_fpregs_23__10_,
         decode_regfile_fpregs_23__11_, decode_regfile_fpregs_23__12_,
         decode_regfile_fpregs_23__13_, decode_regfile_fpregs_23__14_,
         decode_regfile_fpregs_23__15_, decode_regfile_fpregs_23__16_,
         decode_regfile_fpregs_23__17_, decode_regfile_fpregs_23__18_,
         decode_regfile_fpregs_23__19_, decode_regfile_fpregs_23__20_,
         decode_regfile_fpregs_23__21_, decode_regfile_fpregs_23__22_,
         decode_regfile_fpregs_23__23_, decode_regfile_fpregs_23__24_,
         decode_regfile_fpregs_23__25_, decode_regfile_fpregs_23__26_,
         decode_regfile_fpregs_23__27_, decode_regfile_fpregs_23__28_,
         decode_regfile_fpregs_23__29_, decode_regfile_fpregs_23__30_,
         decode_regfile_fpregs_23__31_, decode_regfile_fpregs_24__0_,
         decode_regfile_fpregs_24__1_, decode_regfile_fpregs_24__2_,
         decode_regfile_fpregs_24__3_, decode_regfile_fpregs_24__4_,
         decode_regfile_fpregs_24__5_, decode_regfile_fpregs_24__6_,
         decode_regfile_fpregs_24__7_, decode_regfile_fpregs_24__8_,
         decode_regfile_fpregs_24__9_, decode_regfile_fpregs_24__10_,
         decode_regfile_fpregs_24__11_, decode_regfile_fpregs_24__12_,
         decode_regfile_fpregs_24__13_, decode_regfile_fpregs_24__14_,
         decode_regfile_fpregs_24__15_, decode_regfile_fpregs_24__16_,
         decode_regfile_fpregs_24__17_, decode_regfile_fpregs_24__18_,
         decode_regfile_fpregs_24__19_, decode_regfile_fpregs_24__20_,
         decode_regfile_fpregs_24__21_, decode_regfile_fpregs_24__22_,
         decode_regfile_fpregs_24__23_, decode_regfile_fpregs_24__24_,
         decode_regfile_fpregs_24__25_, decode_regfile_fpregs_24__26_,
         decode_regfile_fpregs_24__27_, decode_regfile_fpregs_24__28_,
         decode_regfile_fpregs_24__29_, decode_regfile_fpregs_24__30_,
         decode_regfile_fpregs_24__31_, decode_regfile_fpregs_25__0_,
         decode_regfile_fpregs_25__1_, decode_regfile_fpregs_25__2_,
         decode_regfile_fpregs_25__3_, decode_regfile_fpregs_25__4_,
         decode_regfile_fpregs_25__5_, decode_regfile_fpregs_25__6_,
         decode_regfile_fpregs_25__7_, decode_regfile_fpregs_25__8_,
         decode_regfile_fpregs_25__9_, decode_regfile_fpregs_25__10_,
         decode_regfile_fpregs_25__11_, decode_regfile_fpregs_25__12_,
         decode_regfile_fpregs_25__13_, decode_regfile_fpregs_25__14_,
         decode_regfile_fpregs_25__15_, decode_regfile_fpregs_25__16_,
         decode_regfile_fpregs_25__17_, decode_regfile_fpregs_25__18_,
         decode_regfile_fpregs_25__19_, decode_regfile_fpregs_25__20_,
         decode_regfile_fpregs_25__21_, decode_regfile_fpregs_25__22_,
         decode_regfile_fpregs_25__23_, decode_regfile_fpregs_25__24_,
         decode_regfile_fpregs_25__25_, decode_regfile_fpregs_25__26_,
         decode_regfile_fpregs_25__27_, decode_regfile_fpregs_25__28_,
         decode_regfile_fpregs_25__29_, decode_regfile_fpregs_25__30_,
         decode_regfile_fpregs_25__31_, decode_regfile_fpregs_26__0_,
         decode_regfile_fpregs_26__1_, decode_regfile_fpregs_26__2_,
         decode_regfile_fpregs_26__3_, decode_regfile_fpregs_26__4_,
         decode_regfile_fpregs_26__5_, decode_regfile_fpregs_26__6_,
         decode_regfile_fpregs_26__7_, decode_regfile_fpregs_26__8_,
         decode_regfile_fpregs_26__9_, decode_regfile_fpregs_26__10_,
         decode_regfile_fpregs_26__11_, decode_regfile_fpregs_26__12_,
         decode_regfile_fpregs_26__13_, decode_regfile_fpregs_26__14_,
         decode_regfile_fpregs_26__15_, decode_regfile_fpregs_26__16_,
         decode_regfile_fpregs_26__17_, decode_regfile_fpregs_26__18_,
         decode_regfile_fpregs_26__19_, decode_regfile_fpregs_26__20_,
         decode_regfile_fpregs_26__21_, decode_regfile_fpregs_26__22_,
         decode_regfile_fpregs_26__23_, decode_regfile_fpregs_26__24_,
         decode_regfile_fpregs_26__25_, decode_regfile_fpregs_26__26_,
         decode_regfile_fpregs_26__27_, decode_regfile_fpregs_26__28_,
         decode_regfile_fpregs_26__29_, decode_regfile_fpregs_26__30_,
         decode_regfile_fpregs_26__31_, decode_regfile_fpregs_27__0_,
         decode_regfile_fpregs_27__1_, decode_regfile_fpregs_27__2_,
         decode_regfile_fpregs_27__3_, decode_regfile_fpregs_27__4_,
         decode_regfile_fpregs_27__5_, decode_regfile_fpregs_27__6_,
         decode_regfile_fpregs_27__7_, decode_regfile_fpregs_27__8_,
         decode_regfile_fpregs_27__9_, decode_regfile_fpregs_27__10_,
         decode_regfile_fpregs_27__11_, decode_regfile_fpregs_27__12_,
         decode_regfile_fpregs_27__13_, decode_regfile_fpregs_27__14_,
         decode_regfile_fpregs_27__15_, decode_regfile_fpregs_27__16_,
         decode_regfile_fpregs_27__17_, decode_regfile_fpregs_27__18_,
         decode_regfile_fpregs_27__19_, decode_regfile_fpregs_27__20_,
         decode_regfile_fpregs_27__21_, decode_regfile_fpregs_27__22_,
         decode_regfile_fpregs_27__23_, decode_regfile_fpregs_27__24_,
         decode_regfile_fpregs_27__25_, decode_regfile_fpregs_27__26_,
         decode_regfile_fpregs_27__27_, decode_regfile_fpregs_27__28_,
         decode_regfile_fpregs_27__29_, decode_regfile_fpregs_27__30_,
         decode_regfile_fpregs_27__31_, decode_regfile_fpregs_28__0_,
         decode_regfile_fpregs_28__1_, decode_regfile_fpregs_28__2_,
         decode_regfile_fpregs_28__3_, decode_regfile_fpregs_28__4_,
         decode_regfile_fpregs_28__5_, decode_regfile_fpregs_28__6_,
         decode_regfile_fpregs_28__7_, decode_regfile_fpregs_28__8_,
         decode_regfile_fpregs_28__9_, decode_regfile_fpregs_28__10_,
         decode_regfile_fpregs_28__11_, decode_regfile_fpregs_28__12_,
         decode_regfile_fpregs_28__13_, decode_regfile_fpregs_28__14_,
         decode_regfile_fpregs_28__15_, decode_regfile_fpregs_28__16_,
         decode_regfile_fpregs_28__17_, decode_regfile_fpregs_28__18_,
         decode_regfile_fpregs_28__19_, decode_regfile_fpregs_28__20_,
         decode_regfile_fpregs_28__21_, decode_regfile_fpregs_28__22_,
         decode_regfile_fpregs_28__23_, decode_regfile_fpregs_28__24_,
         decode_regfile_fpregs_28__25_, decode_regfile_fpregs_28__26_,
         decode_regfile_fpregs_28__27_, decode_regfile_fpregs_28__28_,
         decode_regfile_fpregs_28__29_, decode_regfile_fpregs_28__30_,
         decode_regfile_fpregs_28__31_, decode_regfile_fpregs_29__0_,
         decode_regfile_fpregs_29__1_, decode_regfile_fpregs_29__2_,
         decode_regfile_fpregs_29__3_, decode_regfile_fpregs_29__4_,
         decode_regfile_fpregs_29__5_, decode_regfile_fpregs_29__6_,
         decode_regfile_fpregs_29__7_, decode_regfile_fpregs_29__8_,
         decode_regfile_fpregs_29__9_, decode_regfile_fpregs_29__10_,
         decode_regfile_fpregs_29__11_, decode_regfile_fpregs_29__12_,
         decode_regfile_fpregs_29__13_, decode_regfile_fpregs_29__14_,
         decode_regfile_fpregs_29__15_, decode_regfile_fpregs_29__16_,
         decode_regfile_fpregs_29__17_, decode_regfile_fpregs_29__18_,
         decode_regfile_fpregs_29__19_, decode_regfile_fpregs_29__20_,
         decode_regfile_fpregs_29__21_, decode_regfile_fpregs_29__22_,
         decode_regfile_fpregs_29__23_, decode_regfile_fpregs_29__24_,
         decode_regfile_fpregs_29__25_, decode_regfile_fpregs_29__26_,
         decode_regfile_fpregs_29__27_, decode_regfile_fpregs_29__28_,
         decode_regfile_fpregs_29__29_, decode_regfile_fpregs_29__30_,
         decode_regfile_fpregs_29__31_, decode_regfile_fpregs_30__0_,
         decode_regfile_fpregs_30__1_, decode_regfile_fpregs_30__2_,
         decode_regfile_fpregs_30__3_, decode_regfile_fpregs_30__4_,
         decode_regfile_fpregs_30__5_, decode_regfile_fpregs_30__6_,
         decode_regfile_fpregs_30__7_, decode_regfile_fpregs_30__8_,
         decode_regfile_fpregs_30__9_, decode_regfile_fpregs_30__10_,
         decode_regfile_fpregs_30__11_, decode_regfile_fpregs_30__12_,
         decode_regfile_fpregs_30__13_, decode_regfile_fpregs_30__14_,
         decode_regfile_fpregs_30__15_, decode_regfile_fpregs_30__16_,
         decode_regfile_fpregs_30__17_, decode_regfile_fpregs_30__18_,
         decode_regfile_fpregs_30__19_, decode_regfile_fpregs_30__20_,
         decode_regfile_fpregs_30__21_, decode_regfile_fpregs_30__22_,
         decode_regfile_fpregs_30__23_, decode_regfile_fpregs_30__24_,
         decode_regfile_fpregs_30__25_, decode_regfile_fpregs_30__26_,
         decode_regfile_fpregs_30__27_, decode_regfile_fpregs_30__28_,
         decode_regfile_fpregs_30__29_, decode_regfile_fpregs_30__30_,
         decode_regfile_fpregs_30__31_, decode_regfile_fpregs_31__0_,
         decode_regfile_fpregs_31__1_, decode_regfile_fpregs_31__2_,
         decode_regfile_fpregs_31__3_, decode_regfile_fpregs_31__4_,
         decode_regfile_fpregs_31__5_, decode_regfile_fpregs_31__6_,
         decode_regfile_fpregs_31__7_, decode_regfile_fpregs_31__8_,
         decode_regfile_fpregs_31__9_, decode_regfile_fpregs_31__10_,
         decode_regfile_fpregs_31__11_, decode_regfile_fpregs_31__12_,
         decode_regfile_fpregs_31__13_, decode_regfile_fpregs_31__14_,
         decode_regfile_fpregs_31__15_, decode_regfile_fpregs_31__16_,
         decode_regfile_fpregs_31__17_, decode_regfile_fpregs_31__18_,
         decode_regfile_fpregs_31__19_, decode_regfile_fpregs_31__20_,
         decode_regfile_fpregs_31__21_, decode_regfile_fpregs_31__22_,
         decode_regfile_fpregs_31__23_, decode_regfile_fpregs_31__24_,
         decode_regfile_fpregs_31__25_, decode_regfile_fpregs_31__26_,
         decode_regfile_fpregs_31__27_, decode_regfile_fpregs_31__28_,
         decode_regfile_fpregs_31__29_, decode_regfile_fpregs_31__30_,
         decode_regfile_fpregs_31__31_, execstage_ALUSrc,
         execstage_register_N183, execstage_register_N182,
         execstage_register_N181, execstage_register_N180,
         execstage_register_N179, execstage_register_N178,
         execstage_register_N151, execstage_register_N150,
         execstage_register_N149, execstage_register_N148,
         execstage_register_N147, execstage_register_N146,
         execstage_register_N145, execstage_register_N144,
         execstage_register_N143, execstage_register_N142,
         execstage_register_N141, execstage_register_N140,
         execstage_register_N139, execstage_register_N138,
         execstage_register_N137, execstage_register_N136,
         execstage_register_N135, execstage_register_N134,
         execstage_register_N133, execstage_register_N132,
         execstage_register_N131, execstage_register_N130,
         execstage_register_N129, execstage_register_N128,
         execstage_register_N127, execstage_register_N126,
         execstage_register_N125, execstage_register_N124,
         execstage_register_N123, execstage_register_N122,
         execstage_register_N121, execstage_register_N120,
         execstage_register_N119, execstage_register_N118,
         execstage_register_N117, execstage_register_N116,
         execstage_register_N115, execstage_register_N114,
         execstage_register_N113, execstage_register_N112,
         execstage_register_N111, execstage_register_N110,
         execstage_register_N109, execstage_register_N108,
         execstage_register_N107, execstage_register_N106,
         execstage_register_N105, execstage_register_N104,
         execstage_register_N103, execstage_register_N102,
         execstage_register_N101, execstage_register_N100,
         execstage_register_N99, execstage_register_N98,
         execstage_register_N97, execstage_register_N96,
         execstage_register_N95, execstage_register_N94,
         execstage_register_N93, execstage_register_N92,
         execstage_register_N91, execstage_register_N90,
         execstage_register_N89, execstage_register_N88,
         execstage_register_N87, execstage_register_N86,
         execstage_register_N85, execstage_register_N84,
         execstage_register_N83, execstage_register_N82,
         execstage_register_N81, execstage_register_N80,
         execstage_register_N79, execstage_register_N78,
         execstage_register_N77, execstage_register_N76,
         execstage_register_N75, execstage_register_N74,
         execstage_register_N73, execstage_register_N72,
         execstage_register_N71, execstage_register_N70,
         execstage_register_N69, execstage_register_N68,
         execstage_register_N67, execstage_register_N66,
         execstage_register_N65, execstage_register_N64,
         execstage_register_N63, execstage_register_N62,
         execstage_register_N61, execstage_register_N60,
         execstage_register_N59, execstage_register_N58,
         execstage_register_N57, execstage_register_N56,
         execstage_register_N55, execstage_register_N54,
         execstage_register_N53, execstage_register_N52,
         execstage_register_N51, execstage_register_N50,
         execstage_register_N29, execstage_register_N28,
         execstage_register_N27, execstage_register_N26,
         execstage_register_N25, execstage_register_N23,
         execstage_register_N22, execstage_register_N21,
         execstage_register_N20, execstage_register_N19,
         execstage_register_N18, execstage_register_N14,
         execstage_register_N13, execstage_register_N12,
         execstage_register_N11, execstage_register_N10, execstage_register_N9,
         execstage_register_N6, execstage_register_N5, execstage_register_N4,
         execstage_ALU_N160, execstage_ALU_sel, execstage_ALU_ra_row2_31_,
         mem_memtoreg_out, rgwrite_jalout, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n57, n63, n66, n69, n72, n75, n78, n81, n84, n87,
         n91, n94, n97, n100, n103, n106, n109, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n134, n135, n137, n138, n139, n141,
         n142, n143, n145, n147, n148, n149, n159, n160, n161, n162, n163,
         n191, n202, n215, n220, n222, n225, n228, n231, n234, n237, n240,
         n243, n246, n249, n252, n255, n258, n261, n264, n266, n267, n277,
         n278, n279, n280, n281, n282, n283, n284, n286, n292, n293, n294,
         n296, n299, n300, n301, n302, n304, n305, n306, n309, n312, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n333,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n393,
         n395, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1270, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1471, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2578, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2662, n2663, n2665, n2666, n2667, n2668, n2669, n2672,
         n2673, n2674, n2675, n2677, n2678, n2679, n2681, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2706, n2707, n2708,
         n2710, n2713, n2715, n2717, n2719, n2721, n2723, n2724, n2725, n2726,
         n2727, n2729, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2742, n2743, n2744, n2745, n2746, n2748, n2749, n2750, n2751,
         n2753, n2754, n2755, n2756, n2760, n2762, n2763, n2764, n2765, n2766,
         n2767, n2769, n2770, n2771, n2772, n2773, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2783, n2784, n2785, n2786, n2787, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2799, n2800, n2801, n2802,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2813, n2814,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2825, n2826,
         n2827, n2828, n2830, n2831, n2832, n2833, n2834, n2836, n2837, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2851, n2853, n2854, n2856, n2857, n2858, n2859, n2861, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2872, n2873, n2874, n2878,
         n2880, n2881, n2882, n2883, n2884, n2885, n2887, n2888, n2890, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2900, n2901, n2902, n2903,
         n2906, n2907, n2909, n2911, n2912, n2913, n2915, n2916, n2917, n2919,
         n2920, n2921, n2923, n2924, n2925, n2926, n2927, n2929, n2930, n2931,
         n2932, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2980, n2981, n2982, n2983, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3031, n3032, n3033, n3034, n3036, n3037, n3038, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3103, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3141, n3142, n3143, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3174, n3175, n3176, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3209, n3212, n3213, n3214, n3215, n3216, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3230, n3231, n3232,
         n3234, n3235, n3236, n3237, n3238, n3239, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3259, n3260, n3262, n3263, n3264, n3265, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3275, n3276, n3278, n3279,
         n3281, n3282, n3284, n3285, n3287, n3288, n3290, n3291, n3293, n3294,
         n3295, n3296, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3309, n3310, n3311, n3313, n3314, n3315, n3317, n3318,
         n3319, n3320, n3321, n3323, n3324, n3325, n3326, n3327, n3328, n3330,
         n3331, n3332, n3335, n3336, n3338, n3340, n3341, n3343, n3344, n3345,
         n3347, n3348, n3349, n3351, n3352, n3353, n3355, n3356, n3357, n3360,
         n3361, n3363, n3364, n3365, n3367, n3368, n3370, n3371, n3373, n3374,
         n3375, n3376, n3377, n3379, n3380, n3381, n3382, n3383, n3384, n3386,
         n3387, n3388, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3403, n3404, n3405, n3407, n3408, n3409,
         n3410, n3411, n3412, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3428, n3429, n3430, n3432, n3434, n3435,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3449, n3450, n3451, n3452, n3453, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3467, n3468, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3488, n3489, n3490, n3491, n3492,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3508, n3509, n3510, n3511, n3512, n3513, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3557, n3558,
         n3559, n3560, n3561, n3563, n3564, n3565, n3567, n3568, n3569, n3570,
         n3571, n3573, n3574, n3575, n3576, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3597, n3598, n3599, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3640, n3641, n3643, n3645, n3646, n3647, n3648,
         n3649, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3799, n3801, n3802, n3803,
         n3804, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3945, n3947, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4057, n4058,
         n4059, n4061, n4062, n4063, n4065, n4066, n4068, n4069, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4114, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4137, n4138, n4139,
         n4140, n4142, n4143, n4144, n4145, n4147, n4148, n4149, n4150, n4152,
         n4153, n4154, n4155, n4157, n4158, n4159, n4160, n4162, n4163, n4164,
         n4165, n4167, n4168, n4169, n4170, n4171, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4245, n4246, n4247, n4248, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4261, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4282, n4283, n4284, n4285,
         n4286, n4288, n4289, n4290, n4291, n4292, n4294, n4295, n4296, n4297,
         n4298, n4300, n4301, n4302, n4303, n4304, n4306, n4307, n4308, n4309,
         n4310, n4312, n4313, n4314, n4315, n4316, n4318, n4319, n4320, n4321,
         n4322, n4323, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4423, n4424, n4425, n4426,
         n4427, n4429, n4430, n4431, n4432, n4433, n4435, n4436, n4437, n4438,
         n4439, n4441, n4442, n4443, n4444, n4445, n4447, n4448, n4449, n4450,
         n4451, n4453, n4454, n4455, n4456, n4457, n4459, n4460, n4461, n4462,
         n4463, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4526, n4527, n4529, n4530, n4531, n4532, n4533, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4575, n4576, n4577, n4578, n4579, n4581,
         n4582, n4583, n4584, n4585, n4587, n4588, n4589, n4590, n4591, n4593,
         n4594, n4595, n4596, n4597, n4599, n4600, n4601, n4602, n4603, n4604,
         n4606, n4607, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4627,
         n4628, n4629, n4631, n4632, n4633, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4662, n4664, n4666, n4667, n4668, n4669, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4705,
         n4706, n4707, n4708, n4709, n4711, n4712, n4713, n4714, n4715, n4717,
         n4718, n4719, n4720, n4721, n4723, n4724, n4725, n4726, n4727, n4729,
         n4730, n4731, n4732, n4733, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4755, n4756, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4794,
         n4795, n4796, n4797, n4798, n4799, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4839,
         n4840, n4841, n4842, n4843, n4845, n4846, n4847, n4848, n4849, n4851,
         n4852, n4853, n4854, n4855, n4857, n4858, n4859, n4860, n4861, n4862,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4939, n4940, n4941, n4943, n4944, n4945, n4947, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4983, n4984, n4985, n4986, n4987, n4989, n4990, n4991,
         n4992, n4993, n4995, n4996, n4997, n4998, n4999, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5052, n5054, n5055, n5057,
         n5058, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5107, n5108, n5109, n5110, n5111,
         n5112, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5266, n5267, n5268, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5366, n5367, n5368, n5369, n5371, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5396, n5397,
         n5398, n5399, n5400, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5446, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5458, n5459, n5460, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5484, n5485,
         n5486, n5487, n5488, n5489, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5528, n5529, n5530, n5533, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5587, n5588, n5589, n5590, n5591, n5592,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5611, n5612, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5622, n5625, n5626, n5628, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5650, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5668, n5669, n5670, n5671, n5672, n5673, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5708,
         n5709, n5712, n5715, n5717, n5718, n5719, n5720, n5721, n5722, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5787, n5788,
         n5790, n5791, n5792, n5793, n5795, n5796, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5982,
         n5983, n5984, n5985, n5986, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6017, n6018, n6019, n6020, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6030, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6047, n6049,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6068, n6069, n6070, n6072,
         n6073, n6074, n6076, n6077, n6078, n6079, n6081, n6082, n6084, n6085,
         n6086, n6087, n6088, n6090, n6091, n6093, n6094, n6095, n6096, n6098,
         n6099, n6101, n6102, n6103, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6119, n6120, n6122,
         n6124, n6125, n6126, n6127, n6128, n6129, n6131, n6132, n6133, n6134,
         n6135, n6137, n6138, n6139, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6168, n6169, n6170, n6171, n6172, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6186, n6187, n6188, n6189, n6190, n6191,
         n6193, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n16152, n16153, n16154, n16155, n16156, n16157, n16158,
         n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
         n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174,
         n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182,
         n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190,
         n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198,
         n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206,
         n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214,
         n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222,
         n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230,
         n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238,
         n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246,
         n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254,
         n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262,
         n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270,
         n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278,
         n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286,
         n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294,
         n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302,
         n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
         n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318,
         n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326,
         n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
         n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342,
         n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
         n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358,
         n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366,
         n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374,
         n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
         n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
         n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398,
         n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406,
         n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414,
         n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422,
         n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430,
         n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438,
         n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446,
         n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,
         n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462,
         n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470,
         n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478,
         n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486,
         n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494,
         n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502,
         n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510,
         n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518,
         n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526,
         n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534,
         n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542,
         n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550,
         n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558,
         n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566,
         n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574,
         n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582,
         n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590,
         n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598,
         n16599, n16600, n16601, n16602, n16603, n16604, n16605;
  wire   [4:0] rw_3;
  wire   [1:0] fpoint_3;
  wire   [31:16] instruction_1;
  wire   [15:0] imm32_0;
  wire   [31:0] aluout_0;
  wire   [1:0] fwdA;
  wire   [1:0] fwdB;
  wire   [3:0] aluctrl_0;
  wire   [31:27] instruction_2;
  wire   [4:0] rw_1;
  wire   [1:0] fpoint_1;
  wire   [31:0] busB_1;
  wire   [31:0] delayslot2_2;
  wire   [1:0] fpoint_2;
  wire   [4:0] rw_2;
  wire   [31:0] delayslot2_3;
  wire   [30:0] execstage_BusA;
  wire   [31:0] execstage_Imm32;
  wire   [3:0] execstage_AluCtrl;
  wire   [31:0] mem_ExecResult;
  wire   [31:0] rgwrite_delayslot2out;
  wire   [31:0] rgwrite_busWout;

  AND2_X2 C275 ( .A1(n16371), .A2(N139), .ZN(N38) );
  AND2_X2 C260 ( .A1(n16371), .A2(N139), .ZN(N23) );
  AND2_X2 C248 ( .A1(n13808), .A2(clock), .ZN(N15) );
  OAI33_X1 U5054 ( .A1(n2866), .A2(n13201), .A3(n13227), .B1(n2870), .B2(
        n13188), .B3(n16551), .ZN(n2868) );
  OAI33_X1 U7583 ( .A1(n5642), .A2(n2851), .A3(n13201), .B1(n5547), .B2(n13162), .B3(n13227), .ZN(n5638) );
  OAI33_X1 U8296 ( .A1(n13151), .A2(n13199), .A3(n3418), .B1(n16478), .B2(
        n13102), .B3(n8712), .ZN(n6158) );
  DFF_X2 rgwrite_writereg_qrw_reg_4_ ( .D(rw_2[4]), .CK(clock), .Q(rw_3[4]), 
        .QN(n8753) );
  DFF_X2 execstage_register_qBusB_reg_17_ ( .D(execstage_register_N100), .CK(
        clock), .Q(busB_1[17]) );
  DFF_X2 mem_mRegister_qExecResult_reg_19_ ( .D(aluout_0[19]), .CK(clock), .Q(
        mem_ExecResult[19]) );
  DFF_X2 execstage_register_qRegWrite_reg ( .D(execstage_register_N6), .CK(
        clock), .Q(regwrite_1) );
  DFF_X2 mem_mRegister_qRegWr_reg ( .D(regwrite_1), .CK(clock), .Q(regwrite_2)
         );
  DLH_X2 fwdA_reg_0_ ( .G(N27), .D(n16216), .Q(fwdA[0]) );
  DLH_X2 stall_reg ( .G(N46), .D(N47), .Q(stall) );
  DFF_X2 execstage_register_qMemToReg_reg ( .D(execstage_register_N5), .CK(
        clock), .Q(mem2reg_1) );
  DFF_X2 mem_mRegister_qMemtoReg_reg ( .D(mem2reg_1), .CK(clock), .Q(
        mem_memtoreg_out), .QN(n8725) );
  DFF_X2 rgwrite_writereg_qbusW_reg_19_ ( .D(n16213), .CK(clock), .Q(
        rgwrite_busWout[19]) );
  DFF_X2 execstage_register_qImm32_reg_9_ ( .D(execstage_register_N28), .CK(
        clock), .Q(execstage_Imm32[9]) );
  DFF_X2 execstage_register_qImm32_reg_8_ ( .D(execstage_register_N27), .CK(
        clock), .Q(execstage_Imm32[8]) );
  DFF_X2 execstage_register_qImm32_reg_5_ ( .D(n16218), .CK(clock), .Q(
        execstage_Imm32[5]) );
  DFF_X2 execstage_register_qFPoint_reg_1_ ( .D(execstage_register_N14), .CK(
        clock), .Q(fpoint_1[1]) );
  DFF_X2 mem_mRegister_qFPoint_reg_1_ ( .D(fpoint_1[1]), .CK(clock), .Q(
        fpoint_2[1]) );
  DFF_X2 rgwrite_writereg_qfpoint_reg_1_ ( .D(fpoint_2[1]), .CK(clock), .Q(
        fpoint_3[1]), .QN(n8724) );
  DFF_X2 execstage_register_qFPoint_reg_0_ ( .D(execstage_register_N13), .CK(
        clock), .Q(fpoint_1[0]) );
  DFF_X2 mem_mRegister_qFPoint_reg_0_ ( .D(fpoint_1[0]), .CK(clock), .Q(
        fpoint_2[0]) );
  DFF_X2 rgwrite_writereg_qfpoint_reg_0_ ( .D(fpoint_2[0]), .CK(clock), .Q(
        fpoint_3[0]) );
  DFF_X2 execstage_register_qImm32_reg_15_ ( .D(n16219), .CK(clock), .Q(
        execstage_Imm32[15]) );
  DFF_X2 execstage_register_qImm32_reg_14_ ( .D(n16220), .CK(clock), .Q(
        execstage_Imm32[14]) );
  DFF_X2 execstage_register_qImm32_reg_13_ ( .D(n16221), .CK(clock), .Q(
        execstage_Imm32[13]) );
  DFF_X2 execstage_register_qImm32_reg_12_ ( .D(n16222), .CK(clock), .Q(
        execstage_Imm32[12]) );
  DFF_X2 execstage_register_qRw_reg_4_ ( .D(execstage_register_N119), .CK(
        clock), .Q(rw_1[4]) );
  DFF_X2 mem_mRegister_qRw_reg_4_ ( .D(rw_1[4]), .CK(clock), .Q(rw_2[4]) );
  DFF_X2 execstage_register_qRw_reg_3_ ( .D(execstage_register_N118), .CK(
        clock), .Q(rw_1[3]) );
  DFF_X2 mem_mRegister_qRw_reg_3_ ( .D(rw_1[3]), .CK(clock), .Q(rw_2[3]) );
  DFF_X2 rgwrite_writereg_qrw_reg_3_ ( .D(rw_2[3]), .CK(clock), .Q(rw_3[3]), 
        .QN(n8752) );
  DFF_X2 execstage_register_qRw_reg_2_ ( .D(execstage_register_N117), .CK(
        clock), .Q(rw_1[2]) );
  DFF_X2 mem_mRegister_qRw_reg_2_ ( .D(rw_1[2]), .CK(clock), .Q(rw_2[2]) );
  DFF_X2 rgwrite_writereg_qrw_reg_2_ ( .D(rw_2[2]), .CK(clock), .Q(rw_3[2]), 
        .QN(n8729) );
  DFF_X2 execstage_register_qRw_reg_1_ ( .D(execstage_register_N116), .CK(
        clock), .Q(rw_1[1]), .QN(n8796) );
  DFF_X2 mem_mRegister_qRw_reg_1_ ( .D(rw_1[1]), .CK(clock), .Q(rw_2[1]), .QN(
        n8806) );
  DFF_X2 rgwrite_writereg_qrw_reg_1_ ( .D(rw_2[1]), .CK(clock), .Q(rw_3[1]), 
        .QN(n8755) );
  DFF_X2 execstage_register_qImm32_reg_11_ ( .D(n16223), .CK(clock), .Q(
        execstage_Imm32[11]) );
  DFF_X2 execstage_register_qRw_reg_0_ ( .D(execstage_register_N115), .CK(
        clock), .Q(rw_1[0]), .QN(n8795) );
  DFF_X2 mem_mRegister_qRw_reg_0_ ( .D(rw_1[0]), .CK(clock), .Q(rw_2[0]), .QN(
        n8803) );
  DFF_X2 rgwrite_writereg_qrw_reg_0_ ( .D(rw_2[0]), .CK(clock), .Q(rw_3[0]), 
        .QN(n8754) );
  DLH_X2 stallack_reg ( .G(N14), .D(N15), .Q(stallack) );
  DFF_X2 execstage_register_qBusA_reg_19_ ( .D(execstage_register_N70), .CK(
        clock), .Q(execstage_BusA[19]), .QN(n8654) );
  DFF_X2 execstage_register_qALUSrc_reg ( .D(execstage_register_N4), .CK(clock), .Q(execstage_ALUSrc), .QN(n8708) );
  DFF_X2 execstage_register_qImm32_reg_10_ ( .D(execstage_register_N29), .CK(
        clock), .Q(execstage_Imm32[10]) );
  DFF_X2 execstage_register_qImm32_reg_7_ ( .D(execstage_register_N26), .CK(
        clock), .Q(execstage_Imm32[7]) );
  DFF_X2 execstage_register_qImm32_reg_6_ ( .D(execstage_register_N25), .CK(
        clock), .Q(execstage_Imm32[6]) );
  DFF_X2 execstage_register_qImm32_reg_4_ ( .D(execstage_register_N23), .CK(
        clock), .Q(execstage_Imm32[4]) );
  DFF_X2 execstage_register_qImm32_reg_3_ ( .D(execstage_register_N22), .CK(
        clock), .Q(execstage_Imm32[3]) );
  DFF_X2 execstage_register_qImm32_reg_2_ ( .D(execstage_register_N21), .CK(
        clock), .Q(execstage_Imm32[2]) );
  DFF_X2 execstage_register_qImm32_reg_1_ ( .D(execstage_register_N20), .CK(
        clock), .Q(execstage_Imm32[1]) );
  DFF_X2 execstage_register_qImm32_reg_0_ ( .D(execstage_register_N19), .CK(
        clock), .Q(execstage_Imm32[0]) );
  DFF_X2 execstage_register_qInst_reg_31_ ( .D(execstage_register_N183), .CK(
        clock), .Q(instruction_2[31]) );
  DFF_X2 execstage_register_qInst_reg_30_ ( .D(execstage_register_N182), .CK(
        clock), .Q(instruction_2[30]) );
  DFF_X2 execstage_register_qInst_reg_29_ ( .D(execstage_register_N181), .CK(
        clock), .Q(instruction_2[29]), .QN(n8797) );
  DFF_X2 execstage_register_qInst_reg_28_ ( .D(execstage_register_N180), .CK(
        clock), .Q(instruction_2[28]) );
  DFF_X2 execstage_register_qInst_reg_27_ ( .D(execstage_register_N179), .CK(
        clock), .Q(instruction_2[27]) );
  DFF_X2 execstage_register_qInst_reg_26_ ( .D(execstage_register_N178), .CK(
        clock), .QN(n8762) );
  DLH_X2 fwdB_reg_0_ ( .G(N43), .D(n16215), .Q(fwdB[0]) );
  DLH_X2 fwdB_reg_1_ ( .G(N43), .D(N44), .Q(fwdB[1]) );
  DLH_X2 fwdA_reg_1_ ( .G(N27), .D(N28), .Q(fwdA[1]) );
  DFF_X2 execstage_register_qImm32_reg_31_ ( .D(execstage_register_N50), .CK(
        clock), .Q(execstage_Imm32[31]) );
  DFF_X2 execstage_register_qImm32_reg_29_ ( .D(execstage_register_N50), .CK(
        clock), .Q(execstage_Imm32[29]) );
  DFF_X2 execstage_register_qImm32_reg_27_ ( .D(execstage_register_N50), .CK(
        clock), .Q(execstage_Imm32[27]) );
  DFF_X2 execstage_register_qImm32_reg_25_ ( .D(execstage_register_N50), .CK(
        clock), .Q(execstage_Imm32[25]) );
  DFF_X2 execstage_register_qImm32_reg_23_ ( .D(execstage_register_N50), .CK(
        clock), .Q(execstage_Imm32[23]) );
  DFF_X2 execstage_register_qImm32_reg_21_ ( .D(execstage_register_N50), .CK(
        clock), .Q(execstage_Imm32[21]) );
  DFF_X2 execstage_register_qImm32_reg_19_ ( .D(execstage_register_N50), .CK(
        clock), .Q(execstage_Imm32[19]) );
  DFF_X2 execstage_register_qImm32_reg_17_ ( .D(execstage_register_N50), .CK(
        clock), .Q(execstage_Imm32[17]) );
  DFF_X2 execstage_register_qImm32_reg_16_ ( .D(execstage_register_N50), .CK(
        clock), .Q(execstage_Imm32[16]) );
  DFF_X2 execstage_register_qImm32_reg_18_ ( .D(execstage_register_N50), .CK(
        clock), .Q(execstage_Imm32[18]) );
  DFF_X2 execstage_register_qImm32_reg_20_ ( .D(execstage_register_N50), .CK(
        clock), .Q(execstage_Imm32[20]) );
  DFF_X2 execstage_register_qImm32_reg_22_ ( .D(execstage_register_N50), .CK(
        clock), .Q(execstage_Imm32[22]) );
  DFF_X2 execstage_register_qImm32_reg_24_ ( .D(execstage_register_N50), .CK(
        clock), .Q(execstage_Imm32[24]) );
  DFF_X2 execstage_register_qImm32_reg_26_ ( .D(execstage_register_N50), .CK(
        clock), .Q(execstage_Imm32[26]) );
  DFF_X2 execstage_register_qImm32_reg_28_ ( .D(execstage_register_N50), .CK(
        clock), .Q(execstage_Imm32[28]) );
  DFF_X2 execstage_register_qImm32_reg_30_ ( .D(execstage_register_N50), .CK(
        clock), .Q(execstage_Imm32[30]) );
  DLH_X2 decode_decoder_aluctl_reg_0_ ( .G(decode_decoder_N275), .D(
        decode_decoder_N276), .Q(aluctrl_0[0]) );
  DFF_X2 execstage_register_qAluCtrl_reg_0_ ( .D(execstage_register_N9), .CK(
        clock), .Q(execstage_AluCtrl[0]) );
  DLH_X2 decode_decoder_aluctl_reg_1_ ( .G(decode_decoder_N275), .D(
        decode_decoder_N277), .Q(aluctrl_0[1]) );
  DFF_X2 execstage_register_qAluCtrl_reg_1_ ( .D(execstage_register_N10), .CK(
        clock), .Q(execstage_AluCtrl[1]), .QN(n8720) );
  DLH_X2 decode_decoder_aluctl_reg_2_ ( .G(decode_decoder_N275), .D(
        decode_decoder_N278), .Q(aluctrl_0[2]) );
  DFF_X2 execstage_register_qAluCtrl_reg_2_ ( .D(execstage_register_N11), .CK(
        clock), .Q(execstage_AluCtrl[2]), .QN(n8697) );
  DLH_X2 decode_decoder_aluctl_reg_3_ ( .G(decode_decoder_N275), .D(
        decode_decoder_N279), .Q(aluctrl_0[3]) );
  DFF_X2 execstage_register_qAluCtrl_reg_3_ ( .D(execstage_register_N12), .CK(
        clock), .Q(execstage_AluCtrl[3]), .QN(n8660) );
  DLH_X2 execstage_ALU_sel_reg ( .G(execstage_ALU_N160), .D(n16550), .Q(
        execstage_ALU_sel) );
  DLH_X2 decode_decoder_jall_reg ( .G(decode_decoder_N273), .D(
        decode_decoder_N274), .Q(jal_0) );
  DFF_X2 execstage_register_qJal_reg ( .D(execstage_register_N18), .CK(clock), 
        .Q(jal_1) );
  DFF_X2 mem_mRegister_qJal_reg ( .D(jal_1), .CK(clock), .Q(jal_2) );
  DFF_X2 rgwrite_writereg_qjal_reg ( .D(jal_2), .CK(clock), .Q(rgwrite_jalout), 
        .QN(n8721) );
  DFF_X2 execstage_register_qDelayslot2_reg_0_ ( .D(execstage_register_N120), 
        .CK(clock), .Q(delayslot2_2[0]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_0_ ( .D(delayslot2_2[0]), .CK(clock), 
        .Q(delayslot2_3[0]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_0_ ( .D(delayslot2_3[0]), .CK(clock), 
        .Q(rgwrite_delayslot2out[0]) );
  DFF_X2 execstage_register_qDelayslot2_reg_1_ ( .D(execstage_register_N121), 
        .CK(clock), .Q(delayslot2_2[1]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_1_ ( .D(delayslot2_2[1]), .CK(clock), 
        .Q(delayslot2_3[1]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_1_ ( .D(delayslot2_3[1]), .CK(clock), 
        .Q(rgwrite_delayslot2out[1]) );
  DFF_X2 execstage_register_qDelayslot2_reg_2_ ( .D(execstage_register_N122), 
        .CK(clock), .Q(delayslot2_2[2]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_2_ ( .D(delayslot2_2[2]), .CK(clock), 
        .Q(delayslot2_3[2]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_2_ ( .D(delayslot2_3[2]), .CK(clock), 
        .Q(rgwrite_delayslot2out[2]) );
  DFF_X2 execstage_register_qDelayslot2_reg_3_ ( .D(execstage_register_N123), 
        .CK(clock), .Q(delayslot2_2[3]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_3_ ( .D(delayslot2_2[3]), .CK(clock), 
        .Q(delayslot2_3[3]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_3_ ( .D(delayslot2_3[3]), .CK(clock), 
        .Q(rgwrite_delayslot2out[3]) );
  DFF_X2 execstage_register_qDelayslot2_reg_4_ ( .D(execstage_register_N124), 
        .CK(clock), .Q(delayslot2_2[4]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_4_ ( .D(delayslot2_2[4]), .CK(clock), 
        .Q(delayslot2_3[4]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_4_ ( .D(delayslot2_3[4]), .CK(clock), 
        .Q(rgwrite_delayslot2out[4]) );
  DFF_X2 execstage_register_qDelayslot2_reg_5_ ( .D(execstage_register_N125), 
        .CK(clock), .Q(delayslot2_2[5]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_5_ ( .D(delayslot2_2[5]), .CK(clock), 
        .Q(delayslot2_3[5]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_5_ ( .D(delayslot2_3[5]), .CK(clock), 
        .Q(rgwrite_delayslot2out[5]) );
  DFF_X2 execstage_register_qDelayslot2_reg_6_ ( .D(execstage_register_N126), 
        .CK(clock), .Q(delayslot2_2[6]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_6_ ( .D(delayslot2_2[6]), .CK(clock), 
        .Q(delayslot2_3[6]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_6_ ( .D(delayslot2_3[6]), .CK(clock), 
        .Q(rgwrite_delayslot2out[6]) );
  DFF_X2 execstage_register_qDelayslot2_reg_7_ ( .D(execstage_register_N127), 
        .CK(clock), .Q(delayslot2_2[7]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_7_ ( .D(delayslot2_2[7]), .CK(clock), 
        .Q(delayslot2_3[7]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_7_ ( .D(delayslot2_3[7]), .CK(clock), 
        .Q(rgwrite_delayslot2out[7]) );
  DFF_X2 execstage_register_qDelayslot2_reg_8_ ( .D(execstage_register_N128), 
        .CK(clock), .Q(delayslot2_2[8]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_8_ ( .D(delayslot2_2[8]), .CK(clock), 
        .Q(delayslot2_3[8]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_8_ ( .D(delayslot2_3[8]), .CK(clock), 
        .Q(rgwrite_delayslot2out[8]) );
  DFF_X2 execstage_register_qDelayslot2_reg_9_ ( .D(execstage_register_N129), 
        .CK(clock), .Q(delayslot2_2[9]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_9_ ( .D(delayslot2_2[9]), .CK(clock), 
        .Q(delayslot2_3[9]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_9_ ( .D(delayslot2_3[9]), .CK(clock), 
        .Q(rgwrite_delayslot2out[9]) );
  DFF_X2 execstage_register_qDelayslot2_reg_10_ ( .D(execstage_register_N130), 
        .CK(clock), .Q(delayslot2_2[10]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_10_ ( .D(delayslot2_2[10]), .CK(clock), 
        .Q(delayslot2_3[10]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_10_ ( .D(delayslot2_3[10]), .CK(
        clock), .Q(rgwrite_delayslot2out[10]) );
  DFF_X2 execstage_register_qDelayslot2_reg_11_ ( .D(execstage_register_N131), 
        .CK(clock), .Q(delayslot2_2[11]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_11_ ( .D(delayslot2_2[11]), .CK(clock), 
        .Q(delayslot2_3[11]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_11_ ( .D(delayslot2_3[11]), .CK(
        clock), .Q(rgwrite_delayslot2out[11]) );
  DFF_X2 execstage_register_qDelayslot2_reg_12_ ( .D(execstage_register_N132), 
        .CK(clock), .Q(delayslot2_2[12]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_12_ ( .D(delayslot2_2[12]), .CK(clock), 
        .Q(delayslot2_3[12]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_12_ ( .D(delayslot2_3[12]), .CK(
        clock), .Q(rgwrite_delayslot2out[12]) );
  DFF_X2 execstage_register_qDelayslot2_reg_13_ ( .D(execstage_register_N133), 
        .CK(clock), .Q(delayslot2_2[13]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_13_ ( .D(delayslot2_2[13]), .CK(clock), 
        .Q(delayslot2_3[13]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_13_ ( .D(delayslot2_3[13]), .CK(
        clock), .Q(rgwrite_delayslot2out[13]) );
  DFF_X2 execstage_register_qDelayslot2_reg_14_ ( .D(execstage_register_N134), 
        .CK(clock), .Q(delayslot2_2[14]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_14_ ( .D(delayslot2_2[14]), .CK(clock), 
        .Q(delayslot2_3[14]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_14_ ( .D(delayslot2_3[14]), .CK(
        clock), .Q(rgwrite_delayslot2out[14]) );
  DFF_X2 execstage_register_qDelayslot2_reg_15_ ( .D(execstage_register_N135), 
        .CK(clock), .Q(delayslot2_2[15]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_15_ ( .D(delayslot2_2[15]), .CK(clock), 
        .Q(delayslot2_3[15]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_15_ ( .D(delayslot2_3[15]), .CK(
        clock), .Q(rgwrite_delayslot2out[15]) );
  DFF_X2 execstage_register_qDelayslot2_reg_16_ ( .D(execstage_register_N136), 
        .CK(clock), .Q(delayslot2_2[16]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_16_ ( .D(delayslot2_2[16]), .CK(clock), 
        .Q(delayslot2_3[16]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_16_ ( .D(delayslot2_3[16]), .CK(
        clock), .Q(rgwrite_delayslot2out[16]) );
  DFF_X2 execstage_register_qDelayslot2_reg_17_ ( .D(execstage_register_N137), 
        .CK(clock), .Q(delayslot2_2[17]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_17_ ( .D(delayslot2_2[17]), .CK(clock), 
        .Q(delayslot2_3[17]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_17_ ( .D(delayslot2_3[17]), .CK(
        clock), .Q(rgwrite_delayslot2out[17]) );
  DFF_X2 execstage_register_qDelayslot2_reg_18_ ( .D(execstage_register_N138), 
        .CK(clock), .Q(delayslot2_2[18]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_18_ ( .D(delayslot2_2[18]), .CK(clock), 
        .Q(delayslot2_3[18]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_18_ ( .D(delayslot2_3[18]), .CK(
        clock), .Q(rgwrite_delayslot2out[18]) );
  DFF_X2 execstage_register_qDelayslot2_reg_19_ ( .D(execstage_register_N139), 
        .CK(clock), .Q(delayslot2_2[19]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_19_ ( .D(delayslot2_2[19]), .CK(clock), 
        .Q(delayslot2_3[19]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_19_ ( .D(delayslot2_3[19]), .CK(
        clock), .Q(rgwrite_delayslot2out[19]) );
  DFF_X2 execstage_register_qBusB_reg_19_ ( .D(execstage_register_N102), .CK(
        clock), .Q(busB_1[19]) );
  DFF_X2 execstage_register_qDelayslot2_reg_20_ ( .D(execstage_register_N140), 
        .CK(clock), .Q(delayslot2_2[20]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_20_ ( .D(delayslot2_2[20]), .CK(clock), 
        .Q(delayslot2_3[20]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_20_ ( .D(delayslot2_3[20]), .CK(
        clock), .Q(rgwrite_delayslot2out[20]) );
  DFF_X2 execstage_register_qDelayslot2_reg_21_ ( .D(execstage_register_N141), 
        .CK(clock), .Q(delayslot2_2[21]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_21_ ( .D(delayslot2_2[21]), .CK(clock), 
        .Q(delayslot2_3[21]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_21_ ( .D(delayslot2_3[21]), .CK(
        clock), .Q(rgwrite_delayslot2out[21]) );
  DFF_X2 execstage_register_qDelayslot2_reg_22_ ( .D(execstage_register_N142), 
        .CK(clock), .Q(delayslot2_2[22]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_22_ ( .D(delayslot2_2[22]), .CK(clock), 
        .Q(delayslot2_3[22]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_22_ ( .D(delayslot2_3[22]), .CK(
        clock), .Q(rgwrite_delayslot2out[22]) );
  DFF_X2 execstage_register_qDelayslot2_reg_23_ ( .D(execstage_register_N143), 
        .CK(clock), .Q(delayslot2_2[23]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_23_ ( .D(delayslot2_2[23]), .CK(clock), 
        .Q(delayslot2_3[23]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_23_ ( .D(delayslot2_3[23]), .CK(
        clock), .Q(rgwrite_delayslot2out[23]) );
  DFF_X2 execstage_register_qDelayslot2_reg_24_ ( .D(execstage_register_N144), 
        .CK(clock), .Q(delayslot2_2[24]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_24_ ( .D(delayslot2_2[24]), .CK(clock), 
        .Q(delayslot2_3[24]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_24_ ( .D(delayslot2_3[24]), .CK(
        clock), .Q(rgwrite_delayslot2out[24]) );
  DFF_X2 execstage_register_qDelayslot2_reg_25_ ( .D(execstage_register_N145), 
        .CK(clock), .Q(delayslot2_2[25]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_25_ ( .D(delayslot2_2[25]), .CK(clock), 
        .Q(delayslot2_3[25]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_25_ ( .D(delayslot2_3[25]), .CK(
        clock), .Q(rgwrite_delayslot2out[25]) );
  DFF_X2 execstage_register_qDelayslot2_reg_26_ ( .D(execstage_register_N146), 
        .CK(clock), .Q(delayslot2_2[26]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_26_ ( .D(delayslot2_2[26]), .CK(clock), 
        .Q(delayslot2_3[26]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_26_ ( .D(delayslot2_3[26]), .CK(
        clock), .Q(rgwrite_delayslot2out[26]) );
  DFF_X2 execstage_register_qDelayslot2_reg_27_ ( .D(execstage_register_N147), 
        .CK(clock), .Q(delayslot2_2[27]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_27_ ( .D(delayslot2_2[27]), .CK(clock), 
        .Q(delayslot2_3[27]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_27_ ( .D(delayslot2_3[27]), .CK(
        clock), .Q(rgwrite_delayslot2out[27]) );
  DFF_X2 execstage_register_qDelayslot2_reg_28_ ( .D(execstage_register_N148), 
        .CK(clock), .Q(delayslot2_2[28]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_28_ ( .D(delayslot2_2[28]), .CK(clock), 
        .Q(delayslot2_3[28]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_28_ ( .D(delayslot2_3[28]), .CK(
        clock), .Q(rgwrite_delayslot2out[28]) );
  DFF_X2 execstage_register_qDelayslot2_reg_29_ ( .D(execstage_register_N149), 
        .CK(clock), .Q(delayslot2_2[29]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_29_ ( .D(delayslot2_2[29]), .CK(clock), 
        .Q(delayslot2_3[29]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_29_ ( .D(delayslot2_3[29]), .CK(
        clock), .Q(rgwrite_delayslot2out[29]) );
  DFF_X2 execstage_register_qDelayslot2_reg_30_ ( .D(execstage_register_N150), 
        .CK(clock), .Q(delayslot2_2[30]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_30_ ( .D(delayslot2_2[30]), .CK(clock), 
        .Q(delayslot2_3[30]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_30_ ( .D(delayslot2_3[30]), .CK(
        clock), .Q(rgwrite_delayslot2out[30]) );
  DFF_X2 execstage_register_qDelayslot2_reg_31_ ( .D(execstage_register_N151), 
        .CK(clock), .Q(delayslot2_2[31]) );
  DFF_X2 mem_mRegister_qDelayslot2_reg_31_ ( .D(delayslot2_2[31]), .CK(clock), 
        .Q(delayslot2_3[31]) );
  DFF_X2 rgwrite_writereg_qdelayslot2_reg_31_ ( .D(delayslot2_3[31]), .CK(
        clock), .Q(rgwrite_delayslot2out[31]) );
  DFF_X2 execstage_register_qBusB_reg_31_ ( .D(execstage_register_N114), .CK(
        clock), .Q(busB_1[31]) );
  DFF_X2 mem_mRegister_qExecResult_reg_0_ ( .D(aluout_0[0]), .CK(clock), .Q(
        mem_ExecResult[0]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_0_ ( .D(n16236), .CK(clock), .Q(
        rgwrite_busWout[0]) );
  DFF_X2 execstage_register_qBusB_reg_0_ ( .D(execstage_register_N83), .CK(
        clock), .Q(busB_1[0]) );
  DFF_X2 execstage_register_qBusA_reg_0_ ( .D(execstage_register_N51), .CK(
        clock), .Q(execstage_BusA[0]), .QN(n8712) );
  DFF_X2 mem_mRegister_qExecResult_reg_28_ ( .D(aluout_0[28]), .CK(clock), .Q(
        mem_ExecResult[28]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_28_ ( .D(n16254), .CK(clock), .Q(
        rgwrite_busWout[28]) );
  DFF_X2 execstage_register_qBusB_reg_28_ ( .D(execstage_register_N111), .CK(
        clock), .Q(busB_1[28]) );
  DFF_X2 execstage_register_qBusA_reg_28_ ( .D(execstage_register_N79), .CK(
        clock), .Q(execstage_BusA[28]), .QN(n8735) );
  DFF_X2 mem_mRegister_qExecResult_reg_10_ ( .D(aluout_0[10]), .CK(clock), .Q(
        mem_ExecResult[10]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_10_ ( .D(n16230), .CK(clock), .Q(
        rgwrite_busWout[10]) );
  DFF_X2 execstage_register_qBusB_reg_10_ ( .D(execstage_register_N93), .CK(
        clock), .Q(busB_1[10]) );
  DFF_X2 execstage_register_qBusA_reg_10_ ( .D(execstage_register_N61), .CK(
        clock), .Q(n8694), .QN(n8709) );
  DFF_X2 mem_mRegister_qExecResult_reg_12_ ( .D(aluout_0[12]), .CK(clock), .Q(
        mem_ExecResult[12]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_12_ ( .D(n16224), .CK(clock), .Q(
        rgwrite_busWout[12]) );
  DFF_X2 execstage_register_qBusB_reg_12_ ( .D(execstage_register_N95), .CK(
        clock), .Q(busB_1[12]) );
  DFF_X2 execstage_register_qBusA_reg_12_ ( .D(execstage_register_N63), .CK(
        clock), .Q(execstage_BusA[12]), .QN(n8695) );
  DFF_X2 mem_mRegister_qExecResult_reg_14_ ( .D(aluout_0[14]), .CK(clock), .Q(
        mem_ExecResult[14]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_14_ ( .D(n16226), .CK(clock), .Q(
        rgwrite_busWout[14]) );
  DFF_X2 execstage_register_qBusB_reg_14_ ( .D(execstage_register_N97), .CK(
        clock), .Q(busB_1[14]) );
  DFF_X2 execstage_register_qBusA_reg_14_ ( .D(execstage_register_N65), .CK(
        clock), .Q(execstage_BusA[14]), .QN(n8657) );
  DFF_X2 mem_mRegister_qExecResult_reg_16_ ( .D(aluout_0[16]), .CK(clock), .Q(
        mem_ExecResult[16]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_16_ ( .D(n16244), .CK(clock), .Q(
        rgwrite_busWout[16]) );
  DFF_X2 execstage_register_qBusB_reg_16_ ( .D(execstage_register_N99), .CK(
        clock), .Q(busB_1[16]) );
  DFF_X2 execstage_register_qBusA_reg_16_ ( .D(execstage_register_N67), .CK(
        clock), .Q(execstage_BusA[16]), .QN(n8734) );
  DFF_X2 mem_mRegister_qExecResult_reg_3_ ( .D(aluout_0[3]), .CK(clock), .Q(
        mem_ExecResult[3]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_3_ ( .D(n16239), .CK(clock), .Q(
        rgwrite_busWout[3]) );
  DFF_X2 execstage_register_qBusB_reg_3_ ( .D(execstage_register_N86), .CK(
        clock), .Q(busB_1[3]) );
  DFF_X2 execstage_register_qBusA_reg_3_ ( .D(execstage_register_N54), .CK(
        clock), .Q(n8651), .QN(n8740) );
  DFF_X2 mem_mRegister_qExecResult_reg_4_ ( .D(aluout_0[4]), .CK(clock), .Q(
        mem_ExecResult[4]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_4_ ( .D(n16232), .CK(clock), .Q(
        rgwrite_busWout[4]) );
  DFF_X2 execstage_register_qBusB_reg_4_ ( .D(execstage_register_N87), .CK(
        clock), .Q(busB_1[4]) );
  DFF_X2 execstage_register_qBusA_reg_4_ ( .D(execstage_register_N55), .CK(
        clock), .Q(execstage_BusA[4]), .QN(n8738) );
  DFF_X2 mem_mRegister_qExecResult_reg_11_ ( .D(aluout_0[11]), .CK(clock), .Q(
        mem_ExecResult[11]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_11_ ( .D(n16231), .CK(clock), .Q(
        rgwrite_busWout[11]) );
  DFF_X2 execstage_register_qBusB_reg_11_ ( .D(execstage_register_N94), .CK(
        clock), .Q(busB_1[11]) );
  DFF_X2 execstage_register_qBusA_reg_11_ ( .D(execstage_register_N62), .CK(
        clock), .Q(n8652), .QN(n8736) );
  DFF_X2 mem_mRegister_qExecResult_reg_13_ ( .D(aluout_0[13]), .CK(clock), .Q(
        mem_ExecResult[13]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_13_ ( .D(n16225), .CK(clock), .Q(
        rgwrite_busWout[13]) );
  DFF_X2 execstage_register_qBusB_reg_13_ ( .D(execstage_register_N96), .CK(
        clock), .Q(busB_1[13]) );
  DFF_X2 execstage_register_qBusA_reg_13_ ( .D(execstage_register_N64), .CK(
        clock), .Q(n8655), .QN(n8710) );
  DFF_X2 mem_mRegister_qExecResult_reg_5_ ( .D(aluout_0[5]), .CK(clock), .Q(
        mem_ExecResult[5]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_5_ ( .D(n16233), .CK(clock), .Q(
        rgwrite_busWout[5]) );
  DFF_X2 execstage_register_qBusB_reg_5_ ( .D(execstage_register_N88), .CK(
        clock), .Q(busB_1[5]) );
  DFF_X2 execstage_register_qBusA_reg_5_ ( .D(execstage_register_N56), .CK(
        clock), .Q(execstage_BusA[5]), .QN(n8693) );
  DFF_X2 mem_mRegister_qExecResult_reg_9_ ( .D(aluout_0[9]), .CK(clock), .Q(
        mem_ExecResult[9]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_9_ ( .D(n16229), .CK(clock), .Q(
        rgwrite_busWout[9]) );
  DFF_X2 execstage_register_qBusB_reg_9_ ( .D(execstage_register_N92), .CK(
        clock), .Q(busB_1[9]) );
  DFF_X2 execstage_register_qBusA_reg_9_ ( .D(execstage_register_N60), .CK(
        clock), .Q(n8648), .QN(n8711) );
  DFF_X2 mem_mRegister_qExecResult_reg_15_ ( .D(aluout_0[15]), .CK(clock), .Q(
        mem_ExecResult[15]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_15_ ( .D(n16227), .CK(clock), .Q(
        rgwrite_busWout[15]) );
  DFF_X2 execstage_register_qBusB_reg_15_ ( .D(execstage_register_N98), .CK(
        clock), .Q(busB_1[15]) );
  DFF_X2 execstage_register_qBusA_reg_15_ ( .D(execstage_register_N66), .CK(
        clock), .Q(execstage_BusA[15]), .QN(n8645) );
  DFF_X2 mem_mRegister_qExecResult_reg_17_ ( .D(aluout_0[17]), .CK(clock), .Q(
        mem_ExecResult[17]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_17_ ( .D(n16245), .CK(clock), .Q(
        rgwrite_busWout[17]) );
  DFF_X2 execstage_register_qBusA_reg_17_ ( .D(execstage_register_N68), .CK(
        clock), .Q(execstage_BusA[17]), .QN(n8647) );
  DFF_X2 mem_mRegister_qExecResult_reg_21_ ( .D(aluout_0[21]), .CK(clock), .Q(
        mem_ExecResult[21]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_21_ ( .D(n16243), .CK(clock), .Q(
        rgwrite_busWout[21]) );
  DFF_X2 execstage_register_qBusB_reg_21_ ( .D(execstage_register_N104), .CK(
        clock), .Q(busB_1[21]) );
  DFF_X2 execstage_register_qBusA_reg_21_ ( .D(execstage_register_N72), .CK(
        clock), .Q(execstage_BusA[21]), .QN(n8646) );
  DFF_X2 mem_mRegister_qExecResult_reg_22_ ( .D(aluout_0[22]), .CK(clock), .Q(
        mem_ExecResult[22]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_22_ ( .D(n16241), .CK(clock), .Q(
        rgwrite_busWout[22]) );
  DFF_X2 execstage_register_qBusB_reg_22_ ( .D(execstage_register_N105), .CK(
        clock), .Q(busB_1[22]) );
  DFF_X2 execstage_register_qBusA_reg_22_ ( .D(execstage_register_N73), .CK(
        clock), .Q(execstage_BusA[22]), .QN(n8653) );
  DFF_X2 mem_mRegister_qExecResult_reg_23_ ( .D(aluout_0[23]), .CK(clock), .Q(
        mem_ExecResult[23]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_23_ ( .D(n16240), .CK(clock), .Q(
        rgwrite_busWout[23]) );
  DFF_X2 execstage_register_qBusB_reg_23_ ( .D(execstage_register_N106), .CK(
        clock), .Q(busB_1[23]) );
  DFF_X2 execstage_register_qBusA_reg_23_ ( .D(execstage_register_N74), .CK(
        clock), .Q(execstage_BusA[23]), .QN(n8656) );
  DFF_X2 mem_mRegister_qExecResult_reg_24_ ( .D(aluout_0[24]), .CK(clock), .Q(
        mem_ExecResult[24]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_24_ ( .D(n16250), .CK(clock), .Q(
        rgwrite_busWout[24]) );
  DFF_X2 execstage_register_qBusB_reg_24_ ( .D(execstage_register_N107), .CK(
        clock), .Q(busB_1[24]) );
  DFF_X2 execstage_register_qBusA_reg_24_ ( .D(execstage_register_N75), .CK(
        clock), .Q(execstage_BusA[24]), .QN(n8731) );
  DFF_X2 mem_mRegister_qExecResult_reg_20_ ( .D(aluout_0[20]), .CK(clock), .Q(
        mem_ExecResult[20]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_20_ ( .D(n16242), .CK(clock), .Q(
        rgwrite_busWout[20]) );
  DFF_X2 execstage_register_qBusB_reg_20_ ( .D(execstage_register_N103), .CK(
        clock), .Q(busB_1[20]) );
  DFF_X2 execstage_register_qBusA_reg_20_ ( .D(execstage_register_N71), .CK(
        clock), .Q(execstage_BusA[20]), .QN(n8730) );
  DFF_X2 mem_mRegister_qExecResult_reg_25_ ( .D(aluout_0[25]), .CK(clock), .Q(
        mem_ExecResult[25]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_25_ ( .D(n16249), .CK(clock), .Q(
        rgwrite_busWout[25]) );
  DFF_X2 execstage_register_qBusB_reg_25_ ( .D(execstage_register_N108), .CK(
        clock), .Q(busB_1[25]) );
  DFF_X2 execstage_register_qBusA_reg_25_ ( .D(execstage_register_N76), .CK(
        clock), .Q(execstage_BusA[25]), .QN(n8732) );
  DFF_X2 mem_mRegister_qExecResult_reg_26_ ( .D(aluout_0[26]), .CK(clock), .Q(
        mem_ExecResult[26]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_26_ ( .D(n16248), .CK(clock), .Q(
        rgwrite_busWout[26]) );
  DFF_X2 execstage_register_qBusB_reg_26_ ( .D(execstage_register_N109), .CK(
        clock), .Q(busB_1[26]) );
  DFF_X2 execstage_register_qBusA_reg_26_ ( .D(execstage_register_N77), .CK(
        clock), .Q(execstage_BusA[26]), .QN(n8733) );
  DFF_X2 mem_mRegister_qExecResult_reg_27_ ( .D(aluout_0[27]), .CK(clock), .Q(
        mem_ExecResult[27]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_27_ ( .D(n16247), .CK(clock), .Q(
        rgwrite_busWout[27]) );
  DFF_X2 execstage_register_qBusB_reg_27_ ( .D(execstage_register_N110), .CK(
        clock), .Q(busB_1[27]) );
  DFF_X2 execstage_register_qBusA_reg_27_ ( .D(execstage_register_N78), .CK(
        clock), .Q(execstage_BusA[27]), .QN(n8713) );
  DFF_X2 mem_mRegister_qExecResult_reg_29_ ( .D(aluout_0[29]), .CK(clock), .Q(
        mem_ExecResult[29]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_29_ ( .D(n16253), .CK(clock), .Q(
        rgwrite_busWout[29]) );
  DFF_X2 execstage_register_qBusB_reg_29_ ( .D(execstage_register_N112), .CK(
        clock), .Q(busB_1[29]) );
  DFF_X2 execstage_register_qBusA_reg_29_ ( .D(execstage_register_N80), .CK(
        clock), .Q(execstage_BusA[29]), .QN(n8737) );
  DFF_X2 mem_mRegister_qExecResult_reg_8_ ( .D(aluout_0[8]), .CK(clock), .Q(
        mem_ExecResult[8]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_8_ ( .D(n16228), .CK(clock), .Q(
        rgwrite_busWout[8]) );
  DFF_X2 execstage_register_qBusB_reg_8_ ( .D(execstage_register_N91), .CK(
        clock), .Q(busB_1[8]) );
  DFF_X2 execstage_register_qBusA_reg_8_ ( .D(execstage_register_N59), .CK(
        clock), .Q(execstage_BusA[8]), .QN(n8714) );
  DFF_X2 mem_mRegister_qExecResult_reg_18_ ( .D(aluout_0[18]), .CK(clock), .Q(
        mem_ExecResult[18]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_18_ ( .D(n16246), .CK(clock), .Q(
        rgwrite_busWout[18]) );
  DFF_X2 execstage_register_qBusB_reg_18_ ( .D(execstage_register_N101), .CK(
        clock), .Q(busB_1[18]) );
  DFF_X2 execstage_register_qBusA_reg_18_ ( .D(execstage_register_N69), .CK(
        clock), .Q(execstage_BusA[18]), .QN(n8650) );
  DFF_X2 mem_mRegister_qExecResult_reg_30_ ( .D(aluout_0[30]), .CK(clock), .Q(
        mem_ExecResult[30]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_30_ ( .D(n16252), .CK(clock), .Q(
        rgwrite_busWout[30]) );
  DFF_X2 execstage_register_qBusB_reg_30_ ( .D(execstage_register_N113), .CK(
        clock), .Q(busB_1[30]) );
  DFF_X2 execstage_register_qBusA_reg_30_ ( .D(execstage_register_N81), .CK(
        clock), .Q(execstage_BusA[30]), .QN(n8658) );
  DFF_X2 mem_mRegister_qExecResult_reg_1_ ( .D(aluout_0[1]), .CK(clock), .Q(
        mem_ExecResult[1]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_1_ ( .D(n16237), .CK(clock), .Q(
        rgwrite_busWout[1]) );
  DFF_X2 execstage_register_qBusB_reg_1_ ( .D(execstage_register_N84), .CK(
        clock), .Q(busB_1[1]) );
  DFF_X2 execstage_register_qBusA_reg_1_ ( .D(execstage_register_N52), .CK(
        clock), .Q(execstage_BusA[1]) );
  DFF_X2 mem_mRegister_qExecResult_reg_2_ ( .D(aluout_0[2]), .CK(clock), .Q(
        mem_ExecResult[2]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_2_ ( .D(n16238), .CK(clock), .Q(
        rgwrite_busWout[2]) );
  DFF_X2 execstage_register_qBusB_reg_2_ ( .D(execstage_register_N85), .CK(
        clock), .Q(busB_1[2]) );
  DFF_X2 execstage_register_qBusA_reg_2_ ( .D(execstage_register_N53), .CK(
        clock), .Q(execstage_BusA[2]), .QN(n8692) );
  DFF_X2 mem_mRegister_qExecResult_reg_31_ ( .D(aluout_0[31]), .CK(clock), .Q(
        mem_ExecResult[31]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_31_ ( .D(n16251), .CK(clock), .Q(
        rgwrite_busWout[31]) );
  DFF_X2 execstage_register_qBusA_reg_31_ ( .D(execstage_register_N82), .CK(
        clock), .Q(execstage_ALU_ra_row2_31_), .QN(n8744) );
  DFF_X2 mem_mRegister_qExecResult_reg_6_ ( .D(aluout_0[6]), .CK(clock), .Q(
        mem_ExecResult[6]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_6_ ( .D(n16234), .CK(clock), .Q(
        rgwrite_busWout[6]) );
  DFF_X2 execstage_register_qBusB_reg_6_ ( .D(execstage_register_N89), .CK(
        clock), .Q(busB_1[6]) );
  DFF_X2 execstage_register_qBusA_reg_6_ ( .D(execstage_register_N57), .CK(
        clock), .Q(execstage_BusA[6]), .QN(n8715) );
  DFF_X2 mem_mRegister_qExecResult_reg_7_ ( .D(aluout_0[7]), .CK(clock), .Q(
        mem_ExecResult[7]) );
  DFF_X2 rgwrite_writereg_qbusW_reg_7_ ( .D(n16235), .CK(clock), .Q(
        rgwrite_busWout[7]) );
  DFF_X2 execstage_register_qBusB_reg_7_ ( .D(execstage_register_N90), .CK(
        clock), .Q(busB_1[7]) );
  DFF_X2 execstage_register_qBusA_reg_7_ ( .D(execstage_register_N58), .CK(
        clock), .Q(execstage_BusA[7]), .QN(n8739) );
  DFF_X2 rgwrite_writereg_qregwr_reg ( .D(regwrite_2), .CK(clock), .Q(wrenable) );
  DFF_X2 decode_register_qinst_reg_0_ ( .D(n8306), .CK(clock), .Q(imm32_0[0]), 
        .QN(n8748) );
  DFF_X2 decode_register_qinst_reg_1_ ( .D(n8305), .CK(clock), .Q(imm32_0[1]), 
        .QN(n8726) );
  DFF_X2 decode_register_qinst_reg_2_ ( .D(n8304), .CK(clock), .Q(imm32_0[2]), 
        .QN(n8727) );
  DFF_X2 decode_register_qinst_reg_3_ ( .D(n8303), .CK(clock), .Q(imm32_0[3]), 
        .QN(n8750) );
  DFF_X2 decode_register_qinst_reg_4_ ( .D(n8302), .CK(clock), .Q(imm32_0[4]), 
        .QN(n8749) );
  DFF_X2 decode_register_qinst_reg_5_ ( .D(n8301), .CK(clock), .Q(imm32_0[5]), 
        .QN(n8759) );
  DFF_X2 decode_register_qinst_reg_6_ ( .D(n8300), .CK(clock), .QN(n8751) );
  DFF_X2 decode_register_qinst_reg_7_ ( .D(n8299), .CK(clock), .QN(n8707) );
  DFF_X2 decode_register_qinst_reg_8_ ( .D(n8298), .CK(clock), .Q(imm32_0[8]), 
        .QN(n8761) );
  DFF_X2 decode_register_qinst_reg_9_ ( .D(n8297), .CK(clock), .Q(imm32_0[9]), 
        .QN(n8760) );
  DFF_X2 decode_register_qinst_reg_10_ ( .D(n8296), .CK(clock), .QN(n8728) );
  DFF_X2 decode_register_qinst_reg_11_ ( .D(n8295), .CK(clock), .Q(imm32_0[11]), .QN(n8802) );
  DFF_X2 decode_register_qinst_reg_12_ ( .D(n8294), .CK(clock), .Q(imm32_0[12]), .QN(n8801) );
  DFF_X2 decode_register_qinst_reg_13_ ( .D(n8293), .CK(clock), .Q(imm32_0[13]), .QN(n8800) );
  DFF_X2 decode_register_qinst_reg_14_ ( .D(n8292), .CK(clock), .Q(imm32_0[14]), .QN(n8799) );
  DFF_X2 decode_register_qinst_reg_15_ ( .D(n8291), .CK(clock), .Q(imm32_0[15]), .QN(n8798) );
  DFF_X2 decode_register_qinst_reg_16_ ( .D(n8290), .CK(clock), .Q(
        instruction_1[16]), .QN(n8723) );
  DFF_X2 decode_register_qinst_reg_17_ ( .D(n8289), .CK(clock), .Q(
        instruction_1[17]), .QN(n8804) );
  DFF_X2 decode_register_qinst_reg_18_ ( .D(n8288), .CK(clock), .Q(
        instruction_1[18]), .QN(n8756) );
  DFF_X2 decode_register_qinst_reg_19_ ( .D(n8287), .CK(clock), .Q(
        instruction_1[19]), .QN(n8757) );
  DFF_X2 decode_register_qinst_reg_20_ ( .D(n8286), .CK(clock), .Q(
        instruction_1[20]), .QN(n8758) );
  DFF_X2 decode_register_qinst_reg_21_ ( .D(n8285), .CK(clock), .Q(
        instruction_1[21]), .QN(n8719) );
  DFF_X2 decode_register_qinst_reg_22_ ( .D(n8284), .CK(clock), .Q(
        instruction_1[22]), .QN(n8805) );
  DFF_X2 decode_register_qinst_reg_23_ ( .D(n8283), .CK(clock), .Q(
        instruction_1[23]), .QN(n8745) );
  DFF_X2 decode_register_qinst_reg_24_ ( .D(n8282), .CK(clock), .Q(
        instruction_1[24]), .QN(n8746) );
  DFF_X2 decode_register_qinst_reg_25_ ( .D(n8281), .CK(clock), .Q(
        instruction_1[25]), .QN(n8747) );
  DFF_X2 decode_register_qinst_reg_26_ ( .D(n8280), .CK(clock), .Q(
        instruction_1[26]), .QN(n8716) );
  DFF_X2 decode_register_qinst_reg_27_ ( .D(n8279), .CK(clock), .Q(
        instruction_1[27]), .QN(n8743) );
  DFF_X2 decode_register_qinst_reg_28_ ( .D(n8278), .CK(clock), .Q(
        instruction_1[28]), .QN(n8717) );
  DFF_X2 decode_register_qinst_reg_29_ ( .D(n8277), .CK(clock), .Q(
        instruction_1[29]), .QN(n8742) );
  DFF_X2 decode_register_qinst_reg_30_ ( .D(n8276), .CK(clock), .Q(
        instruction_1[30]), .QN(n8741) );
  DFF_X2 decode_register_qinst_reg_31_ ( .D(n8275), .CK(clock), .Q(
        instruction_1[31]), .QN(n8718) );
  DFF_X2 decode_register_qdelay2_reg_0_ ( .D(n8274), .CK(clock), .QN(n8794) );
  DFF_X2 decode_register_qdelay2_reg_1_ ( .D(n8273), .CK(clock), .QN(n8793) );
  DFF_X2 decode_register_qdelay2_reg_2_ ( .D(n8272), .CK(clock), .QN(n8792) );
  DFF_X2 decode_register_qdelay2_reg_3_ ( .D(n8271), .CK(clock), .QN(n8791) );
  DFF_X2 decode_register_qdelay2_reg_4_ ( .D(n8270), .CK(clock), .QN(n8790) );
  DFF_X2 decode_register_qdelay2_reg_5_ ( .D(n8269), .CK(clock), .QN(n8789) );
  DFF_X2 decode_register_qdelay2_reg_6_ ( .D(n8268), .CK(clock), .QN(n8788) );
  DFF_X2 decode_register_qdelay2_reg_7_ ( .D(n8267), .CK(clock), .QN(n8787) );
  DFF_X2 decode_register_qdelay2_reg_8_ ( .D(n8266), .CK(clock), .QN(n8786) );
  DFF_X2 decode_register_qdelay2_reg_9_ ( .D(n8265), .CK(clock), .QN(n8785) );
  DFF_X2 decode_register_qdelay2_reg_10_ ( .D(n8264), .CK(clock), .QN(n8784)
         );
  DFF_X2 decode_register_qdelay2_reg_11_ ( .D(n8263), .CK(clock), .QN(n8783)
         );
  DFF_X2 decode_register_qdelay2_reg_12_ ( .D(n8262), .CK(clock), .QN(n8782)
         );
  DFF_X2 decode_register_qdelay2_reg_13_ ( .D(n8261), .CK(clock), .QN(n8781)
         );
  DFF_X2 decode_register_qdelay2_reg_14_ ( .D(n8260), .CK(clock), .QN(n8780)
         );
  DFF_X2 decode_register_qdelay2_reg_15_ ( .D(n8259), .CK(clock), .QN(n8779)
         );
  DFF_X2 decode_register_qdelay2_reg_16_ ( .D(n8258), .CK(clock), .QN(n8778)
         );
  DFF_X2 decode_register_qdelay2_reg_17_ ( .D(n8257), .CK(clock), .QN(n8777)
         );
  DFF_X2 decode_register_qdelay2_reg_18_ ( .D(n8256), .CK(clock), .QN(n8776)
         );
  DFF_X2 decode_register_qdelay2_reg_19_ ( .D(n8255), .CK(clock), .QN(n8775)
         );
  DFF_X2 decode_register_qdelay2_reg_20_ ( .D(n8254), .CK(clock), .QN(n8774)
         );
  DFF_X2 decode_register_qdelay2_reg_21_ ( .D(n8253), .CK(clock), .QN(n8773)
         );
  DFF_X2 decode_register_qdelay2_reg_22_ ( .D(n8252), .CK(clock), .QN(n8772)
         );
  DFF_X2 decode_register_qdelay2_reg_23_ ( .D(n8251), .CK(clock), .QN(n8771)
         );
  DFF_X2 decode_register_qdelay2_reg_24_ ( .D(n8250), .CK(clock), .QN(n8770)
         );
  DFF_X2 decode_register_qdelay2_reg_25_ ( .D(n8249), .CK(clock), .QN(n8769)
         );
  DFF_X2 decode_register_qdelay2_reg_26_ ( .D(n8248), .CK(clock), .QN(n8768)
         );
  DFF_X2 decode_register_qdelay2_reg_27_ ( .D(n8247), .CK(clock), .QN(n8767)
         );
  DFF_X2 decode_register_qdelay2_reg_28_ ( .D(n8246), .CK(clock), .QN(n8766)
         );
  DFF_X2 decode_register_qdelay2_reg_29_ ( .D(n8245), .CK(clock), .QN(n8765)
         );
  DFF_X2 decode_register_qdelay2_reg_30_ ( .D(n8244), .CK(clock), .QN(n8764)
         );
  DFF_X2 decode_register_qdelay2_reg_31_ ( .D(n8243), .CK(clock), .QN(n8763)
         );
  DFF_X2 decode_regfile_fpregs_reg_31__0_ ( .D(n8242), .CK(clock), .Q(
        decode_regfile_fpregs_31__0_) );
  DFF_X2 decode_regfile_fpregs_reg_31__1_ ( .D(n8241), .CK(clock), .Q(
        decode_regfile_fpregs_31__1_) );
  DFF_X2 decode_regfile_fpregs_reg_31__2_ ( .D(n8240), .CK(clock), .Q(
        decode_regfile_fpregs_31__2_) );
  DFF_X2 decode_regfile_fpregs_reg_31__3_ ( .D(n8239), .CK(clock), .Q(
        decode_regfile_fpregs_31__3_) );
  DFF_X2 decode_regfile_fpregs_reg_31__4_ ( .D(n8238), .CK(clock), .Q(
        decode_regfile_fpregs_31__4_) );
  DFF_X2 decode_regfile_fpregs_reg_31__5_ ( .D(n8237), .CK(clock), .Q(
        decode_regfile_fpregs_31__5_) );
  DFF_X2 decode_regfile_fpregs_reg_31__6_ ( .D(n8236), .CK(clock), .Q(
        decode_regfile_fpregs_31__6_) );
  DFF_X2 decode_regfile_fpregs_reg_31__7_ ( .D(n8235), .CK(clock), .Q(
        decode_regfile_fpregs_31__7_) );
  DFF_X2 decode_regfile_fpregs_reg_31__8_ ( .D(n8234), .CK(clock), .Q(
        decode_regfile_fpregs_31__8_) );
  DFF_X2 decode_regfile_fpregs_reg_31__9_ ( .D(n8233), .CK(clock), .Q(
        decode_regfile_fpregs_31__9_) );
  DFF_X2 decode_regfile_fpregs_reg_31__10_ ( .D(n8232), .CK(clock), .Q(
        decode_regfile_fpregs_31__10_) );
  DFF_X2 decode_regfile_fpregs_reg_31__11_ ( .D(n8231), .CK(clock), .Q(
        decode_regfile_fpregs_31__11_) );
  DFF_X2 decode_regfile_fpregs_reg_31__12_ ( .D(n8230), .CK(clock), .Q(
        decode_regfile_fpregs_31__12_) );
  DFF_X2 decode_regfile_fpregs_reg_31__13_ ( .D(n8229), .CK(clock), .Q(
        decode_regfile_fpregs_31__13_) );
  DFF_X2 decode_regfile_fpregs_reg_31__14_ ( .D(n8228), .CK(clock), .Q(
        decode_regfile_fpregs_31__14_) );
  DFF_X2 decode_regfile_fpregs_reg_31__15_ ( .D(n8227), .CK(clock), .Q(
        decode_regfile_fpregs_31__15_) );
  DFF_X2 decode_regfile_fpregs_reg_31__16_ ( .D(n8226), .CK(clock), .Q(
        decode_regfile_fpregs_31__16_) );
  DFF_X2 decode_regfile_fpregs_reg_31__17_ ( .D(n8225), .CK(clock), .Q(
        decode_regfile_fpregs_31__17_) );
  DFF_X2 decode_regfile_fpregs_reg_31__18_ ( .D(n8224), .CK(clock), .Q(
        decode_regfile_fpregs_31__18_) );
  DFF_X2 decode_regfile_fpregs_reg_31__19_ ( .D(n8223), .CK(clock), .Q(
        decode_regfile_fpregs_31__19_) );
  DFF_X2 decode_regfile_fpregs_reg_31__20_ ( .D(n8222), .CK(clock), .Q(
        decode_regfile_fpregs_31__20_) );
  DFF_X2 decode_regfile_fpregs_reg_31__21_ ( .D(n8221), .CK(clock), .Q(
        decode_regfile_fpregs_31__21_) );
  DFF_X2 decode_regfile_fpregs_reg_31__22_ ( .D(n8220), .CK(clock), .Q(
        decode_regfile_fpregs_31__22_) );
  DFF_X2 decode_regfile_fpregs_reg_31__23_ ( .D(n8219), .CK(clock), .Q(
        decode_regfile_fpregs_31__23_) );
  DFF_X2 decode_regfile_fpregs_reg_31__24_ ( .D(n8218), .CK(clock), .Q(
        decode_regfile_fpregs_31__24_) );
  DFF_X2 decode_regfile_fpregs_reg_31__25_ ( .D(n8217), .CK(clock), .Q(
        decode_regfile_fpregs_31__25_) );
  DFF_X2 decode_regfile_fpregs_reg_31__26_ ( .D(n8216), .CK(clock), .Q(
        decode_regfile_fpregs_31__26_) );
  DFF_X2 decode_regfile_fpregs_reg_31__27_ ( .D(n8215), .CK(clock), .Q(
        decode_regfile_fpregs_31__27_) );
  DFF_X2 decode_regfile_fpregs_reg_31__28_ ( .D(n8214), .CK(clock), .Q(
        decode_regfile_fpregs_31__28_) );
  DFF_X2 decode_regfile_fpregs_reg_31__29_ ( .D(n8213), .CK(clock), .Q(
        decode_regfile_fpregs_31__29_) );
  DFF_X2 decode_regfile_fpregs_reg_31__30_ ( .D(n8212), .CK(clock), .Q(
        decode_regfile_fpregs_31__30_) );
  DFF_X2 decode_regfile_fpregs_reg_31__31_ ( .D(n8211), .CK(clock), .Q(
        decode_regfile_fpregs_31__31_) );
  DFF_X2 decode_regfile_fpregs_reg_30__0_ ( .D(n8210), .CK(clock), .Q(
        decode_regfile_fpregs_30__0_) );
  DFF_X2 decode_regfile_fpregs_reg_30__1_ ( .D(n8209), .CK(clock), .Q(
        decode_regfile_fpregs_30__1_) );
  DFF_X2 decode_regfile_fpregs_reg_30__2_ ( .D(n8208), .CK(clock), .Q(
        decode_regfile_fpregs_30__2_) );
  DFF_X2 decode_regfile_fpregs_reg_30__3_ ( .D(n8207), .CK(clock), .Q(
        decode_regfile_fpregs_30__3_) );
  DFF_X2 decode_regfile_fpregs_reg_30__4_ ( .D(n8206), .CK(clock), .Q(
        decode_regfile_fpregs_30__4_) );
  DFF_X2 decode_regfile_fpregs_reg_30__5_ ( .D(n8205), .CK(clock), .Q(
        decode_regfile_fpregs_30__5_) );
  DFF_X2 decode_regfile_fpregs_reg_30__6_ ( .D(n8204), .CK(clock), .Q(
        decode_regfile_fpregs_30__6_) );
  DFF_X2 decode_regfile_fpregs_reg_30__7_ ( .D(n8203), .CK(clock), .Q(
        decode_regfile_fpregs_30__7_) );
  DFF_X2 decode_regfile_fpregs_reg_30__8_ ( .D(n8202), .CK(clock), .Q(
        decode_regfile_fpregs_30__8_) );
  DFF_X2 decode_regfile_fpregs_reg_30__9_ ( .D(n8201), .CK(clock), .Q(
        decode_regfile_fpregs_30__9_) );
  DFF_X2 decode_regfile_fpregs_reg_30__10_ ( .D(n8200), .CK(clock), .Q(
        decode_regfile_fpregs_30__10_) );
  DFF_X2 decode_regfile_fpregs_reg_30__11_ ( .D(n8199), .CK(clock), .Q(
        decode_regfile_fpregs_30__11_) );
  DFF_X2 decode_regfile_fpregs_reg_30__12_ ( .D(n8198), .CK(clock), .Q(
        decode_regfile_fpregs_30__12_) );
  DFF_X2 decode_regfile_fpregs_reg_30__13_ ( .D(n8197), .CK(clock), .Q(
        decode_regfile_fpregs_30__13_) );
  DFF_X2 decode_regfile_fpregs_reg_30__14_ ( .D(n8196), .CK(clock), .Q(
        decode_regfile_fpregs_30__14_) );
  DFF_X2 decode_regfile_fpregs_reg_30__15_ ( .D(n8195), .CK(clock), .Q(
        decode_regfile_fpregs_30__15_) );
  DFF_X2 decode_regfile_fpregs_reg_30__16_ ( .D(n8194), .CK(clock), .Q(
        decode_regfile_fpregs_30__16_) );
  DFF_X2 decode_regfile_fpregs_reg_30__17_ ( .D(n8193), .CK(clock), .Q(
        decode_regfile_fpregs_30__17_) );
  DFF_X2 decode_regfile_fpregs_reg_30__18_ ( .D(n8192), .CK(clock), .Q(
        decode_regfile_fpregs_30__18_) );
  DFF_X2 decode_regfile_fpregs_reg_30__19_ ( .D(n8191), .CK(clock), .Q(
        decode_regfile_fpregs_30__19_) );
  DFF_X2 decode_regfile_fpregs_reg_30__20_ ( .D(n8190), .CK(clock), .Q(
        decode_regfile_fpregs_30__20_) );
  DFF_X2 decode_regfile_fpregs_reg_30__21_ ( .D(n8189), .CK(clock), .Q(
        decode_regfile_fpregs_30__21_) );
  DFF_X2 decode_regfile_fpregs_reg_30__22_ ( .D(n8188), .CK(clock), .Q(
        decode_regfile_fpregs_30__22_) );
  DFF_X2 decode_regfile_fpregs_reg_30__23_ ( .D(n8187), .CK(clock), .Q(
        decode_regfile_fpregs_30__23_) );
  DFF_X2 decode_regfile_fpregs_reg_30__24_ ( .D(n8186), .CK(clock), .Q(
        decode_regfile_fpregs_30__24_) );
  DFF_X2 decode_regfile_fpregs_reg_30__25_ ( .D(n8185), .CK(clock), .Q(
        decode_regfile_fpregs_30__25_) );
  DFF_X2 decode_regfile_fpregs_reg_30__26_ ( .D(n8184), .CK(clock), .Q(
        decode_regfile_fpregs_30__26_) );
  DFF_X2 decode_regfile_fpregs_reg_30__27_ ( .D(n8183), .CK(clock), .Q(
        decode_regfile_fpregs_30__27_) );
  DFF_X2 decode_regfile_fpregs_reg_30__28_ ( .D(n8182), .CK(clock), .Q(
        decode_regfile_fpregs_30__28_) );
  DFF_X2 decode_regfile_fpregs_reg_30__29_ ( .D(n8181), .CK(clock), .Q(
        decode_regfile_fpregs_30__29_) );
  DFF_X2 decode_regfile_fpregs_reg_30__30_ ( .D(n8180), .CK(clock), .Q(
        decode_regfile_fpregs_30__30_) );
  DFF_X2 decode_regfile_fpregs_reg_30__31_ ( .D(n8179), .CK(clock), .Q(
        decode_regfile_fpregs_30__31_) );
  DFF_X2 decode_regfile_fpregs_reg_29__0_ ( .D(n8178), .CK(clock), .Q(
        decode_regfile_fpregs_29__0_) );
  DFF_X2 decode_regfile_fpregs_reg_29__1_ ( .D(n8177), .CK(clock), .Q(
        decode_regfile_fpregs_29__1_) );
  DFF_X2 decode_regfile_fpregs_reg_29__2_ ( .D(n8176), .CK(clock), .Q(
        decode_regfile_fpregs_29__2_) );
  DFF_X2 decode_regfile_fpregs_reg_29__3_ ( .D(n8175), .CK(clock), .Q(
        decode_regfile_fpregs_29__3_) );
  DFF_X2 decode_regfile_fpregs_reg_29__4_ ( .D(n8174), .CK(clock), .Q(
        decode_regfile_fpregs_29__4_) );
  DFF_X2 decode_regfile_fpregs_reg_29__5_ ( .D(n8173), .CK(clock), .Q(
        decode_regfile_fpregs_29__5_) );
  DFF_X2 decode_regfile_fpregs_reg_29__6_ ( .D(n8172), .CK(clock), .Q(
        decode_regfile_fpregs_29__6_) );
  DFF_X2 decode_regfile_fpregs_reg_29__7_ ( .D(n8171), .CK(clock), .Q(
        decode_regfile_fpregs_29__7_) );
  DFF_X2 decode_regfile_fpregs_reg_29__8_ ( .D(n8170), .CK(clock), .Q(
        decode_regfile_fpregs_29__8_) );
  DFF_X2 decode_regfile_fpregs_reg_29__9_ ( .D(n8169), .CK(clock), .Q(
        decode_regfile_fpregs_29__9_) );
  DFF_X2 decode_regfile_fpregs_reg_29__10_ ( .D(n8168), .CK(clock), .Q(
        decode_regfile_fpregs_29__10_) );
  DFF_X2 decode_regfile_fpregs_reg_29__11_ ( .D(n8167), .CK(clock), .Q(
        decode_regfile_fpregs_29__11_) );
  DFF_X2 decode_regfile_fpregs_reg_29__12_ ( .D(n8166), .CK(clock), .Q(
        decode_regfile_fpregs_29__12_) );
  DFF_X2 decode_regfile_fpregs_reg_29__13_ ( .D(n8165), .CK(clock), .Q(
        decode_regfile_fpregs_29__13_) );
  DFF_X2 decode_regfile_fpregs_reg_29__14_ ( .D(n8164), .CK(clock), .Q(
        decode_regfile_fpregs_29__14_) );
  DFF_X2 decode_regfile_fpregs_reg_29__15_ ( .D(n8163), .CK(clock), .Q(
        decode_regfile_fpregs_29__15_) );
  DFF_X2 decode_regfile_fpregs_reg_29__16_ ( .D(n8162), .CK(clock), .Q(
        decode_regfile_fpregs_29__16_) );
  DFF_X2 decode_regfile_fpregs_reg_29__17_ ( .D(n8161), .CK(clock), .Q(
        decode_regfile_fpregs_29__17_) );
  DFF_X2 decode_regfile_fpregs_reg_29__18_ ( .D(n8160), .CK(clock), .Q(
        decode_regfile_fpregs_29__18_) );
  DFF_X2 decode_regfile_fpregs_reg_29__19_ ( .D(n8159), .CK(clock), .Q(
        decode_regfile_fpregs_29__19_) );
  DFF_X2 decode_regfile_fpregs_reg_29__20_ ( .D(n8158), .CK(clock), .Q(
        decode_regfile_fpregs_29__20_) );
  DFF_X2 decode_regfile_fpregs_reg_29__21_ ( .D(n8157), .CK(clock), .Q(
        decode_regfile_fpregs_29__21_) );
  DFF_X2 decode_regfile_fpregs_reg_29__22_ ( .D(n8156), .CK(clock), .Q(
        decode_regfile_fpregs_29__22_) );
  DFF_X2 decode_regfile_fpregs_reg_29__23_ ( .D(n8155), .CK(clock), .Q(
        decode_regfile_fpregs_29__23_) );
  DFF_X2 decode_regfile_fpregs_reg_29__24_ ( .D(n8154), .CK(clock), .Q(
        decode_regfile_fpregs_29__24_) );
  DFF_X2 decode_regfile_fpregs_reg_29__25_ ( .D(n8153), .CK(clock), .Q(
        decode_regfile_fpregs_29__25_) );
  DFF_X2 decode_regfile_fpregs_reg_29__26_ ( .D(n8152), .CK(clock), .Q(
        decode_regfile_fpregs_29__26_) );
  DFF_X2 decode_regfile_fpregs_reg_29__27_ ( .D(n8151), .CK(clock), .Q(
        decode_regfile_fpregs_29__27_) );
  DFF_X2 decode_regfile_fpregs_reg_29__28_ ( .D(n8150), .CK(clock), .Q(
        decode_regfile_fpregs_29__28_) );
  DFF_X2 decode_regfile_fpregs_reg_29__29_ ( .D(n8149), .CK(clock), .Q(
        decode_regfile_fpregs_29__29_) );
  DFF_X2 decode_regfile_fpregs_reg_29__30_ ( .D(n8148), .CK(clock), .Q(
        decode_regfile_fpregs_29__30_) );
  DFF_X2 decode_regfile_fpregs_reg_29__31_ ( .D(n8147), .CK(clock), .Q(
        decode_regfile_fpregs_29__31_) );
  DFF_X2 decode_regfile_fpregs_reg_28__0_ ( .D(n8146), .CK(clock), .Q(
        decode_regfile_fpregs_28__0_) );
  DFF_X2 decode_regfile_fpregs_reg_28__1_ ( .D(n8145), .CK(clock), .Q(
        decode_regfile_fpregs_28__1_) );
  DFF_X2 decode_regfile_fpregs_reg_28__2_ ( .D(n8144), .CK(clock), .Q(
        decode_regfile_fpregs_28__2_) );
  DFF_X2 decode_regfile_fpregs_reg_28__3_ ( .D(n8143), .CK(clock), .Q(
        decode_regfile_fpregs_28__3_) );
  DFF_X2 decode_regfile_fpregs_reg_28__4_ ( .D(n8142), .CK(clock), .Q(
        decode_regfile_fpregs_28__4_) );
  DFF_X2 decode_regfile_fpregs_reg_28__5_ ( .D(n8141), .CK(clock), .Q(
        decode_regfile_fpregs_28__5_) );
  DFF_X2 decode_regfile_fpregs_reg_28__6_ ( .D(n8140), .CK(clock), .Q(
        decode_regfile_fpregs_28__6_) );
  DFF_X2 decode_regfile_fpregs_reg_28__7_ ( .D(n8139), .CK(clock), .Q(
        decode_regfile_fpregs_28__7_) );
  DFF_X2 decode_regfile_fpregs_reg_28__8_ ( .D(n8138), .CK(clock), .Q(
        decode_regfile_fpregs_28__8_) );
  DFF_X2 decode_regfile_fpregs_reg_28__9_ ( .D(n8137), .CK(clock), .Q(
        decode_regfile_fpregs_28__9_) );
  DFF_X2 decode_regfile_fpregs_reg_28__10_ ( .D(n8136), .CK(clock), .Q(
        decode_regfile_fpregs_28__10_) );
  DFF_X2 decode_regfile_fpregs_reg_28__11_ ( .D(n8135), .CK(clock), .Q(
        decode_regfile_fpregs_28__11_) );
  DFF_X2 decode_regfile_fpregs_reg_28__12_ ( .D(n8134), .CK(clock), .Q(
        decode_regfile_fpregs_28__12_) );
  DFF_X2 decode_regfile_fpregs_reg_28__13_ ( .D(n8133), .CK(clock), .Q(
        decode_regfile_fpregs_28__13_) );
  DFF_X2 decode_regfile_fpregs_reg_28__14_ ( .D(n8132), .CK(clock), .Q(
        decode_regfile_fpregs_28__14_) );
  DFF_X2 decode_regfile_fpregs_reg_28__15_ ( .D(n8131), .CK(clock), .Q(
        decode_regfile_fpregs_28__15_) );
  DFF_X2 decode_regfile_fpregs_reg_28__16_ ( .D(n8130), .CK(clock), .Q(
        decode_regfile_fpregs_28__16_) );
  DFF_X2 decode_regfile_fpregs_reg_28__17_ ( .D(n8129), .CK(clock), .Q(
        decode_regfile_fpregs_28__17_) );
  DFF_X2 decode_regfile_fpregs_reg_28__18_ ( .D(n8128), .CK(clock), .Q(
        decode_regfile_fpregs_28__18_) );
  DFF_X2 decode_regfile_fpregs_reg_28__19_ ( .D(n8127), .CK(clock), .Q(
        decode_regfile_fpregs_28__19_) );
  DFF_X2 decode_regfile_fpregs_reg_28__20_ ( .D(n8126), .CK(clock), .Q(
        decode_regfile_fpregs_28__20_) );
  DFF_X2 decode_regfile_fpregs_reg_28__21_ ( .D(n8125), .CK(clock), .Q(
        decode_regfile_fpregs_28__21_) );
  DFF_X2 decode_regfile_fpregs_reg_28__22_ ( .D(n8124), .CK(clock), .Q(
        decode_regfile_fpregs_28__22_) );
  DFF_X2 decode_regfile_fpregs_reg_28__23_ ( .D(n8123), .CK(clock), .Q(
        decode_regfile_fpregs_28__23_) );
  DFF_X2 decode_regfile_fpregs_reg_28__24_ ( .D(n8122), .CK(clock), .Q(
        decode_regfile_fpregs_28__24_) );
  DFF_X2 decode_regfile_fpregs_reg_28__25_ ( .D(n8121), .CK(clock), .Q(
        decode_regfile_fpregs_28__25_) );
  DFF_X2 decode_regfile_fpregs_reg_28__26_ ( .D(n8120), .CK(clock), .Q(
        decode_regfile_fpregs_28__26_) );
  DFF_X2 decode_regfile_fpregs_reg_28__27_ ( .D(n8119), .CK(clock), .Q(
        decode_regfile_fpregs_28__27_) );
  DFF_X2 decode_regfile_fpregs_reg_28__28_ ( .D(n8118), .CK(clock), .Q(
        decode_regfile_fpregs_28__28_) );
  DFF_X2 decode_regfile_fpregs_reg_28__29_ ( .D(n8117), .CK(clock), .Q(
        decode_regfile_fpregs_28__29_) );
  DFF_X2 decode_regfile_fpregs_reg_28__30_ ( .D(n8116), .CK(clock), .Q(
        decode_regfile_fpregs_28__30_) );
  DFF_X2 decode_regfile_fpregs_reg_28__31_ ( .D(n8115), .CK(clock), .Q(
        decode_regfile_fpregs_28__31_) );
  DFF_X2 decode_regfile_fpregs_reg_27__0_ ( .D(n8114), .CK(clock), .Q(
        decode_regfile_fpregs_27__0_) );
  DFF_X2 decode_regfile_fpregs_reg_27__1_ ( .D(n8113), .CK(clock), .Q(
        decode_regfile_fpregs_27__1_) );
  DFF_X2 decode_regfile_fpregs_reg_27__2_ ( .D(n8112), .CK(clock), .Q(
        decode_regfile_fpregs_27__2_) );
  DFF_X2 decode_regfile_fpregs_reg_27__3_ ( .D(n8111), .CK(clock), .Q(
        decode_regfile_fpregs_27__3_) );
  DFF_X2 decode_regfile_fpregs_reg_27__4_ ( .D(n8110), .CK(clock), .Q(
        decode_regfile_fpregs_27__4_) );
  DFF_X2 decode_regfile_fpregs_reg_27__5_ ( .D(n8109), .CK(clock), .Q(
        decode_regfile_fpregs_27__5_) );
  DFF_X2 decode_regfile_fpregs_reg_27__6_ ( .D(n8108), .CK(clock), .Q(
        decode_regfile_fpregs_27__6_) );
  DFF_X2 decode_regfile_fpregs_reg_27__7_ ( .D(n8107), .CK(clock), .Q(
        decode_regfile_fpregs_27__7_) );
  DFF_X2 decode_regfile_fpregs_reg_27__8_ ( .D(n8106), .CK(clock), .Q(
        decode_regfile_fpregs_27__8_) );
  DFF_X2 decode_regfile_fpregs_reg_27__9_ ( .D(n8105), .CK(clock), .Q(
        decode_regfile_fpregs_27__9_) );
  DFF_X2 decode_regfile_fpregs_reg_27__10_ ( .D(n8104), .CK(clock), .Q(
        decode_regfile_fpregs_27__10_) );
  DFF_X2 decode_regfile_fpregs_reg_27__11_ ( .D(n8103), .CK(clock), .Q(
        decode_regfile_fpregs_27__11_) );
  DFF_X2 decode_regfile_fpregs_reg_27__12_ ( .D(n8102), .CK(clock), .Q(
        decode_regfile_fpregs_27__12_) );
  DFF_X2 decode_regfile_fpregs_reg_27__13_ ( .D(n8101), .CK(clock), .Q(
        decode_regfile_fpregs_27__13_) );
  DFF_X2 decode_regfile_fpregs_reg_27__14_ ( .D(n8100), .CK(clock), .Q(
        decode_regfile_fpregs_27__14_) );
  DFF_X2 decode_regfile_fpregs_reg_27__15_ ( .D(n8099), .CK(clock), .Q(
        decode_regfile_fpregs_27__15_) );
  DFF_X2 decode_regfile_fpregs_reg_27__16_ ( .D(n8098), .CK(clock), .Q(
        decode_regfile_fpregs_27__16_) );
  DFF_X2 decode_regfile_fpregs_reg_27__17_ ( .D(n8097), .CK(clock), .Q(
        decode_regfile_fpregs_27__17_) );
  DFF_X2 decode_regfile_fpregs_reg_27__18_ ( .D(n8096), .CK(clock), .Q(
        decode_regfile_fpregs_27__18_) );
  DFF_X2 decode_regfile_fpregs_reg_27__19_ ( .D(n8095), .CK(clock), .Q(
        decode_regfile_fpregs_27__19_) );
  DFF_X2 decode_regfile_fpregs_reg_27__20_ ( .D(n8094), .CK(clock), .Q(
        decode_regfile_fpregs_27__20_) );
  DFF_X2 decode_regfile_fpregs_reg_27__21_ ( .D(n8093), .CK(clock), .Q(
        decode_regfile_fpregs_27__21_) );
  DFF_X2 decode_regfile_fpregs_reg_27__22_ ( .D(n8092), .CK(clock), .Q(
        decode_regfile_fpregs_27__22_) );
  DFF_X2 decode_regfile_fpregs_reg_27__23_ ( .D(n8091), .CK(clock), .Q(
        decode_regfile_fpregs_27__23_) );
  DFF_X2 decode_regfile_fpregs_reg_27__24_ ( .D(n8090), .CK(clock), .Q(
        decode_regfile_fpregs_27__24_) );
  DFF_X2 decode_regfile_fpregs_reg_27__25_ ( .D(n8089), .CK(clock), .Q(
        decode_regfile_fpregs_27__25_) );
  DFF_X2 decode_regfile_fpregs_reg_27__26_ ( .D(n8088), .CK(clock), .Q(
        decode_regfile_fpregs_27__26_) );
  DFF_X2 decode_regfile_fpregs_reg_27__27_ ( .D(n8087), .CK(clock), .Q(
        decode_regfile_fpregs_27__27_) );
  DFF_X2 decode_regfile_fpregs_reg_27__28_ ( .D(n8086), .CK(clock), .Q(
        decode_regfile_fpregs_27__28_) );
  DFF_X2 decode_regfile_fpregs_reg_27__29_ ( .D(n8085), .CK(clock), .Q(
        decode_regfile_fpregs_27__29_) );
  DFF_X2 decode_regfile_fpregs_reg_27__30_ ( .D(n8084), .CK(clock), .Q(
        decode_regfile_fpregs_27__30_) );
  DFF_X2 decode_regfile_fpregs_reg_27__31_ ( .D(n8083), .CK(clock), .Q(
        decode_regfile_fpregs_27__31_) );
  DFF_X2 decode_regfile_fpregs_reg_26__0_ ( .D(n8082), .CK(clock), .Q(
        decode_regfile_fpregs_26__0_) );
  DFF_X2 decode_regfile_fpregs_reg_26__1_ ( .D(n8081), .CK(clock), .Q(
        decode_regfile_fpregs_26__1_) );
  DFF_X2 decode_regfile_fpregs_reg_26__2_ ( .D(n8080), .CK(clock), .Q(
        decode_regfile_fpregs_26__2_) );
  DFF_X2 decode_regfile_fpregs_reg_26__3_ ( .D(n8079), .CK(clock), .Q(
        decode_regfile_fpregs_26__3_) );
  DFF_X2 decode_regfile_fpregs_reg_26__4_ ( .D(n8078), .CK(clock), .Q(
        decode_regfile_fpregs_26__4_) );
  DFF_X2 decode_regfile_fpregs_reg_26__5_ ( .D(n8077), .CK(clock), .Q(
        decode_regfile_fpregs_26__5_) );
  DFF_X2 decode_regfile_fpregs_reg_26__6_ ( .D(n8076), .CK(clock), .Q(
        decode_regfile_fpregs_26__6_) );
  DFF_X2 decode_regfile_fpregs_reg_26__7_ ( .D(n8075), .CK(clock), .Q(
        decode_regfile_fpregs_26__7_) );
  DFF_X2 decode_regfile_fpregs_reg_26__8_ ( .D(n8074), .CK(clock), .Q(
        decode_regfile_fpregs_26__8_) );
  DFF_X2 decode_regfile_fpregs_reg_26__9_ ( .D(n8073), .CK(clock), .Q(
        decode_regfile_fpregs_26__9_) );
  DFF_X2 decode_regfile_fpregs_reg_26__10_ ( .D(n8072), .CK(clock), .Q(
        decode_regfile_fpregs_26__10_) );
  DFF_X2 decode_regfile_fpregs_reg_26__11_ ( .D(n8071), .CK(clock), .Q(
        decode_regfile_fpregs_26__11_) );
  DFF_X2 decode_regfile_fpregs_reg_26__12_ ( .D(n8070), .CK(clock), .Q(
        decode_regfile_fpregs_26__12_) );
  DFF_X2 decode_regfile_fpregs_reg_26__13_ ( .D(n8069), .CK(clock), .Q(
        decode_regfile_fpregs_26__13_) );
  DFF_X2 decode_regfile_fpregs_reg_26__14_ ( .D(n8068), .CK(clock), .Q(
        decode_regfile_fpregs_26__14_) );
  DFF_X2 decode_regfile_fpregs_reg_26__15_ ( .D(n8067), .CK(clock), .Q(
        decode_regfile_fpregs_26__15_) );
  DFF_X2 decode_regfile_fpregs_reg_26__16_ ( .D(n8066), .CK(clock), .Q(
        decode_regfile_fpregs_26__16_) );
  DFF_X2 decode_regfile_fpregs_reg_26__17_ ( .D(n8065), .CK(clock), .Q(
        decode_regfile_fpregs_26__17_) );
  DFF_X2 decode_regfile_fpregs_reg_26__18_ ( .D(n8064), .CK(clock), .Q(
        decode_regfile_fpregs_26__18_) );
  DFF_X2 decode_regfile_fpregs_reg_26__19_ ( .D(n8063), .CK(clock), .Q(
        decode_regfile_fpregs_26__19_) );
  DFF_X2 decode_regfile_fpregs_reg_26__20_ ( .D(n8062), .CK(clock), .Q(
        decode_regfile_fpregs_26__20_) );
  DFF_X2 decode_regfile_fpregs_reg_26__21_ ( .D(n8061), .CK(clock), .Q(
        decode_regfile_fpregs_26__21_) );
  DFF_X2 decode_regfile_fpregs_reg_26__22_ ( .D(n8060), .CK(clock), .Q(
        decode_regfile_fpregs_26__22_) );
  DFF_X2 decode_regfile_fpregs_reg_26__23_ ( .D(n8059), .CK(clock), .Q(
        decode_regfile_fpregs_26__23_) );
  DFF_X2 decode_regfile_fpregs_reg_26__24_ ( .D(n8058), .CK(clock), .Q(
        decode_regfile_fpregs_26__24_) );
  DFF_X2 decode_regfile_fpregs_reg_26__25_ ( .D(n8057), .CK(clock), .Q(
        decode_regfile_fpregs_26__25_) );
  DFF_X2 decode_regfile_fpregs_reg_26__26_ ( .D(n8056), .CK(clock), .Q(
        decode_regfile_fpregs_26__26_) );
  DFF_X2 decode_regfile_fpregs_reg_26__27_ ( .D(n8055), .CK(clock), .Q(
        decode_regfile_fpregs_26__27_) );
  DFF_X2 decode_regfile_fpregs_reg_26__28_ ( .D(n8054), .CK(clock), .Q(
        decode_regfile_fpregs_26__28_) );
  DFF_X2 decode_regfile_fpregs_reg_26__29_ ( .D(n8053), .CK(clock), .Q(
        decode_regfile_fpregs_26__29_) );
  DFF_X2 decode_regfile_fpregs_reg_26__30_ ( .D(n8052), .CK(clock), .Q(
        decode_regfile_fpregs_26__30_) );
  DFF_X2 decode_regfile_fpregs_reg_26__31_ ( .D(n8051), .CK(clock), .Q(
        decode_regfile_fpregs_26__31_) );
  DFF_X2 decode_regfile_fpregs_reg_25__0_ ( .D(n8050), .CK(clock), .Q(
        decode_regfile_fpregs_25__0_) );
  DFF_X2 decode_regfile_fpregs_reg_25__1_ ( .D(n8049), .CK(clock), .Q(
        decode_regfile_fpregs_25__1_) );
  DFF_X2 decode_regfile_fpregs_reg_25__2_ ( .D(n8048), .CK(clock), .Q(
        decode_regfile_fpregs_25__2_) );
  DFF_X2 decode_regfile_fpregs_reg_25__3_ ( .D(n8047), .CK(clock), .Q(
        decode_regfile_fpregs_25__3_) );
  DFF_X2 decode_regfile_fpregs_reg_25__4_ ( .D(n8046), .CK(clock), .Q(
        decode_regfile_fpregs_25__4_) );
  DFF_X2 decode_regfile_fpregs_reg_25__5_ ( .D(n8045), .CK(clock), .Q(
        decode_regfile_fpregs_25__5_) );
  DFF_X2 decode_regfile_fpregs_reg_25__6_ ( .D(n8044), .CK(clock), .Q(
        decode_regfile_fpregs_25__6_) );
  DFF_X2 decode_regfile_fpregs_reg_25__7_ ( .D(n8043), .CK(clock), .Q(
        decode_regfile_fpregs_25__7_) );
  DFF_X2 decode_regfile_fpregs_reg_25__8_ ( .D(n8042), .CK(clock), .Q(
        decode_regfile_fpregs_25__8_) );
  DFF_X2 decode_regfile_fpregs_reg_25__9_ ( .D(n8041), .CK(clock), .Q(
        decode_regfile_fpregs_25__9_) );
  DFF_X2 decode_regfile_fpregs_reg_25__10_ ( .D(n8040), .CK(clock), .Q(
        decode_regfile_fpregs_25__10_) );
  DFF_X2 decode_regfile_fpregs_reg_25__11_ ( .D(n8039), .CK(clock), .Q(
        decode_regfile_fpregs_25__11_) );
  DFF_X2 decode_regfile_fpregs_reg_25__12_ ( .D(n8038), .CK(clock), .Q(
        decode_regfile_fpregs_25__12_) );
  DFF_X2 decode_regfile_fpregs_reg_25__13_ ( .D(n8037), .CK(clock), .Q(
        decode_regfile_fpregs_25__13_) );
  DFF_X2 decode_regfile_fpregs_reg_25__14_ ( .D(n8036), .CK(clock), .Q(
        decode_regfile_fpregs_25__14_) );
  DFF_X2 decode_regfile_fpregs_reg_25__15_ ( .D(n8035), .CK(clock), .Q(
        decode_regfile_fpregs_25__15_) );
  DFF_X2 decode_regfile_fpregs_reg_25__16_ ( .D(n8034), .CK(clock), .Q(
        decode_regfile_fpregs_25__16_) );
  DFF_X2 decode_regfile_fpregs_reg_25__17_ ( .D(n8033), .CK(clock), .Q(
        decode_regfile_fpregs_25__17_) );
  DFF_X2 decode_regfile_fpregs_reg_25__18_ ( .D(n8032), .CK(clock), .Q(
        decode_regfile_fpregs_25__18_) );
  DFF_X2 decode_regfile_fpregs_reg_25__19_ ( .D(n8031), .CK(clock), .Q(
        decode_regfile_fpregs_25__19_) );
  DFF_X2 decode_regfile_fpregs_reg_25__20_ ( .D(n8030), .CK(clock), .Q(
        decode_regfile_fpregs_25__20_) );
  DFF_X2 decode_regfile_fpregs_reg_25__21_ ( .D(n8029), .CK(clock), .Q(
        decode_regfile_fpregs_25__21_) );
  DFF_X2 decode_regfile_fpregs_reg_25__22_ ( .D(n8028), .CK(clock), .Q(
        decode_regfile_fpregs_25__22_) );
  DFF_X2 decode_regfile_fpregs_reg_25__23_ ( .D(n8027), .CK(clock), .Q(
        decode_regfile_fpregs_25__23_) );
  DFF_X2 decode_regfile_fpregs_reg_25__24_ ( .D(n8026), .CK(clock), .Q(
        decode_regfile_fpregs_25__24_) );
  DFF_X2 decode_regfile_fpregs_reg_25__25_ ( .D(n8025), .CK(clock), .Q(
        decode_regfile_fpregs_25__25_) );
  DFF_X2 decode_regfile_fpregs_reg_25__26_ ( .D(n8024), .CK(clock), .Q(
        decode_regfile_fpregs_25__26_) );
  DFF_X2 decode_regfile_fpregs_reg_25__27_ ( .D(n8023), .CK(clock), .Q(
        decode_regfile_fpregs_25__27_) );
  DFF_X2 decode_regfile_fpregs_reg_25__28_ ( .D(n8022), .CK(clock), .Q(
        decode_regfile_fpregs_25__28_) );
  DFF_X2 decode_regfile_fpregs_reg_25__29_ ( .D(n8021), .CK(clock), .Q(
        decode_regfile_fpregs_25__29_) );
  DFF_X2 decode_regfile_fpregs_reg_25__30_ ( .D(n8020), .CK(clock), .Q(
        decode_regfile_fpregs_25__30_) );
  DFF_X2 decode_regfile_fpregs_reg_25__31_ ( .D(n8019), .CK(clock), .Q(
        decode_regfile_fpregs_25__31_) );
  DFF_X2 decode_regfile_fpregs_reg_24__0_ ( .D(n8018), .CK(clock), .Q(
        decode_regfile_fpregs_24__0_) );
  DFF_X2 decode_regfile_fpregs_reg_24__1_ ( .D(n8017), .CK(clock), .Q(
        decode_regfile_fpregs_24__1_) );
  DFF_X2 decode_regfile_fpregs_reg_24__2_ ( .D(n8016), .CK(clock), .Q(
        decode_regfile_fpregs_24__2_) );
  DFF_X2 decode_regfile_fpregs_reg_24__3_ ( .D(n8015), .CK(clock), .Q(
        decode_regfile_fpregs_24__3_) );
  DFF_X2 decode_regfile_fpregs_reg_24__4_ ( .D(n8014), .CK(clock), .Q(
        decode_regfile_fpregs_24__4_) );
  DFF_X2 decode_regfile_fpregs_reg_24__5_ ( .D(n8013), .CK(clock), .Q(
        decode_regfile_fpregs_24__5_) );
  DFF_X2 decode_regfile_fpregs_reg_24__6_ ( .D(n8012), .CK(clock), .Q(
        decode_regfile_fpregs_24__6_) );
  DFF_X2 decode_regfile_fpregs_reg_24__7_ ( .D(n8011), .CK(clock), .Q(
        decode_regfile_fpregs_24__7_) );
  DFF_X2 decode_regfile_fpregs_reg_24__8_ ( .D(n8010), .CK(clock), .Q(
        decode_regfile_fpregs_24__8_) );
  DFF_X2 decode_regfile_fpregs_reg_24__9_ ( .D(n8009), .CK(clock), .Q(
        decode_regfile_fpregs_24__9_) );
  DFF_X2 decode_regfile_fpregs_reg_24__10_ ( .D(n8008), .CK(clock), .Q(
        decode_regfile_fpregs_24__10_) );
  DFF_X2 decode_regfile_fpregs_reg_24__11_ ( .D(n8007), .CK(clock), .Q(
        decode_regfile_fpregs_24__11_) );
  DFF_X2 decode_regfile_fpregs_reg_24__12_ ( .D(n8006), .CK(clock), .Q(
        decode_regfile_fpregs_24__12_) );
  DFF_X2 decode_regfile_fpregs_reg_24__13_ ( .D(n8005), .CK(clock), .Q(
        decode_regfile_fpregs_24__13_) );
  DFF_X2 decode_regfile_fpregs_reg_24__14_ ( .D(n8004), .CK(clock), .Q(
        decode_regfile_fpregs_24__14_) );
  DFF_X2 decode_regfile_fpregs_reg_24__15_ ( .D(n8003), .CK(clock), .Q(
        decode_regfile_fpregs_24__15_) );
  DFF_X2 decode_regfile_fpregs_reg_24__16_ ( .D(n8002), .CK(clock), .Q(
        decode_regfile_fpregs_24__16_) );
  DFF_X2 decode_regfile_fpregs_reg_24__17_ ( .D(n8001), .CK(clock), .Q(
        decode_regfile_fpregs_24__17_) );
  DFF_X2 decode_regfile_fpregs_reg_24__18_ ( .D(n8000), .CK(clock), .Q(
        decode_regfile_fpregs_24__18_) );
  DFF_X2 decode_regfile_fpregs_reg_24__19_ ( .D(n7999), .CK(clock), .Q(
        decode_regfile_fpregs_24__19_) );
  DFF_X2 decode_regfile_fpregs_reg_24__20_ ( .D(n7998), .CK(clock), .Q(
        decode_regfile_fpregs_24__20_) );
  DFF_X2 decode_regfile_fpregs_reg_24__21_ ( .D(n7997), .CK(clock), .Q(
        decode_regfile_fpregs_24__21_) );
  DFF_X2 decode_regfile_fpregs_reg_24__22_ ( .D(n7996), .CK(clock), .Q(
        decode_regfile_fpregs_24__22_) );
  DFF_X2 decode_regfile_fpregs_reg_24__23_ ( .D(n7995), .CK(clock), .Q(
        decode_regfile_fpregs_24__23_) );
  DFF_X2 decode_regfile_fpregs_reg_24__24_ ( .D(n7994), .CK(clock), .Q(
        decode_regfile_fpregs_24__24_) );
  DFF_X2 decode_regfile_fpregs_reg_24__25_ ( .D(n7993), .CK(clock), .Q(
        decode_regfile_fpregs_24__25_) );
  DFF_X2 decode_regfile_fpregs_reg_24__26_ ( .D(n7992), .CK(clock), .Q(
        decode_regfile_fpregs_24__26_) );
  DFF_X2 decode_regfile_fpregs_reg_24__27_ ( .D(n7991), .CK(clock), .Q(
        decode_regfile_fpregs_24__27_) );
  DFF_X2 decode_regfile_fpregs_reg_24__28_ ( .D(n7990), .CK(clock), .Q(
        decode_regfile_fpregs_24__28_) );
  DFF_X2 decode_regfile_fpregs_reg_24__29_ ( .D(n7989), .CK(clock), .Q(
        decode_regfile_fpregs_24__29_) );
  DFF_X2 decode_regfile_fpregs_reg_24__30_ ( .D(n7988), .CK(clock), .Q(
        decode_regfile_fpregs_24__30_) );
  DFF_X2 decode_regfile_fpregs_reg_24__31_ ( .D(n7987), .CK(clock), .Q(
        decode_regfile_fpregs_24__31_) );
  DFF_X2 decode_regfile_fpregs_reg_23__0_ ( .D(n7986), .CK(clock), .Q(
        decode_regfile_fpregs_23__0_) );
  DFF_X2 decode_regfile_fpregs_reg_23__1_ ( .D(n7985), .CK(clock), .Q(
        decode_regfile_fpregs_23__1_) );
  DFF_X2 decode_regfile_fpregs_reg_23__2_ ( .D(n7984), .CK(clock), .Q(
        decode_regfile_fpregs_23__2_) );
  DFF_X2 decode_regfile_fpregs_reg_23__3_ ( .D(n7983), .CK(clock), .Q(
        decode_regfile_fpregs_23__3_) );
  DFF_X2 decode_regfile_fpregs_reg_23__4_ ( .D(n7982), .CK(clock), .Q(
        decode_regfile_fpregs_23__4_) );
  DFF_X2 decode_regfile_fpregs_reg_23__5_ ( .D(n7981), .CK(clock), .Q(
        decode_regfile_fpregs_23__5_) );
  DFF_X2 decode_regfile_fpregs_reg_23__6_ ( .D(n7980), .CK(clock), .Q(
        decode_regfile_fpregs_23__6_) );
  DFF_X2 decode_regfile_fpregs_reg_23__7_ ( .D(n7979), .CK(clock), .Q(
        decode_regfile_fpregs_23__7_) );
  DFF_X2 decode_regfile_fpregs_reg_23__8_ ( .D(n7978), .CK(clock), .Q(
        decode_regfile_fpregs_23__8_) );
  DFF_X2 decode_regfile_fpregs_reg_23__9_ ( .D(n7977), .CK(clock), .Q(
        decode_regfile_fpregs_23__9_) );
  DFF_X2 decode_regfile_fpregs_reg_23__10_ ( .D(n7976), .CK(clock), .Q(
        decode_regfile_fpregs_23__10_) );
  DFF_X2 decode_regfile_fpregs_reg_23__11_ ( .D(n7975), .CK(clock), .Q(
        decode_regfile_fpregs_23__11_) );
  DFF_X2 decode_regfile_fpregs_reg_23__12_ ( .D(n7974), .CK(clock), .Q(
        decode_regfile_fpregs_23__12_) );
  DFF_X2 decode_regfile_fpregs_reg_23__13_ ( .D(n7973), .CK(clock), .Q(
        decode_regfile_fpregs_23__13_) );
  DFF_X2 decode_regfile_fpregs_reg_23__14_ ( .D(n7972), .CK(clock), .Q(
        decode_regfile_fpregs_23__14_) );
  DFF_X2 decode_regfile_fpregs_reg_23__15_ ( .D(n7971), .CK(clock), .Q(
        decode_regfile_fpregs_23__15_) );
  DFF_X2 decode_regfile_fpregs_reg_23__16_ ( .D(n7970), .CK(clock), .Q(
        decode_regfile_fpregs_23__16_) );
  DFF_X2 decode_regfile_fpregs_reg_23__17_ ( .D(n7969), .CK(clock), .Q(
        decode_regfile_fpregs_23__17_) );
  DFF_X2 decode_regfile_fpregs_reg_23__18_ ( .D(n7968), .CK(clock), .Q(
        decode_regfile_fpregs_23__18_) );
  DFF_X2 decode_regfile_fpregs_reg_23__19_ ( .D(n7967), .CK(clock), .Q(
        decode_regfile_fpregs_23__19_) );
  DFF_X2 decode_regfile_fpregs_reg_23__20_ ( .D(n7966), .CK(clock), .Q(
        decode_regfile_fpregs_23__20_) );
  DFF_X2 decode_regfile_fpregs_reg_23__21_ ( .D(n7965), .CK(clock), .Q(
        decode_regfile_fpregs_23__21_) );
  DFF_X2 decode_regfile_fpregs_reg_23__22_ ( .D(n7964), .CK(clock), .Q(
        decode_regfile_fpregs_23__22_) );
  DFF_X2 decode_regfile_fpregs_reg_23__23_ ( .D(n7963), .CK(clock), .Q(
        decode_regfile_fpregs_23__23_) );
  DFF_X2 decode_regfile_fpregs_reg_23__24_ ( .D(n7962), .CK(clock), .Q(
        decode_regfile_fpregs_23__24_) );
  DFF_X2 decode_regfile_fpregs_reg_23__25_ ( .D(n7961), .CK(clock), .Q(
        decode_regfile_fpregs_23__25_) );
  DFF_X2 decode_regfile_fpregs_reg_23__26_ ( .D(n7960), .CK(clock), .Q(
        decode_regfile_fpregs_23__26_) );
  DFF_X2 decode_regfile_fpregs_reg_23__27_ ( .D(n7959), .CK(clock), .Q(
        decode_regfile_fpregs_23__27_) );
  DFF_X2 decode_regfile_fpregs_reg_23__28_ ( .D(n7958), .CK(clock), .Q(
        decode_regfile_fpregs_23__28_) );
  DFF_X2 decode_regfile_fpregs_reg_23__29_ ( .D(n7957), .CK(clock), .Q(
        decode_regfile_fpregs_23__29_) );
  DFF_X2 decode_regfile_fpregs_reg_23__30_ ( .D(n7956), .CK(clock), .Q(
        decode_regfile_fpregs_23__30_) );
  DFF_X2 decode_regfile_fpregs_reg_23__31_ ( .D(n7955), .CK(clock), .Q(
        decode_regfile_fpregs_23__31_) );
  DFF_X2 decode_regfile_fpregs_reg_22__0_ ( .D(n7954), .CK(clock), .Q(
        decode_regfile_fpregs_22__0_) );
  DFF_X2 decode_regfile_fpregs_reg_22__1_ ( .D(n7953), .CK(clock), .Q(
        decode_regfile_fpregs_22__1_) );
  DFF_X2 decode_regfile_fpregs_reg_22__2_ ( .D(n7952), .CK(clock), .Q(
        decode_regfile_fpregs_22__2_) );
  DFF_X2 decode_regfile_fpregs_reg_22__3_ ( .D(n7951), .CK(clock), .Q(
        decode_regfile_fpregs_22__3_) );
  DFF_X2 decode_regfile_fpregs_reg_22__4_ ( .D(n7950), .CK(clock), .Q(
        decode_regfile_fpregs_22__4_) );
  DFF_X2 decode_regfile_fpregs_reg_22__5_ ( .D(n7949), .CK(clock), .Q(
        decode_regfile_fpregs_22__5_) );
  DFF_X2 decode_regfile_fpregs_reg_22__6_ ( .D(n7948), .CK(clock), .Q(
        decode_regfile_fpregs_22__6_) );
  DFF_X2 decode_regfile_fpregs_reg_22__7_ ( .D(n7947), .CK(clock), .Q(
        decode_regfile_fpregs_22__7_) );
  DFF_X2 decode_regfile_fpregs_reg_22__8_ ( .D(n7946), .CK(clock), .Q(
        decode_regfile_fpregs_22__8_) );
  DFF_X2 decode_regfile_fpregs_reg_22__9_ ( .D(n7945), .CK(clock), .Q(
        decode_regfile_fpregs_22__9_) );
  DFF_X2 decode_regfile_fpregs_reg_22__10_ ( .D(n7944), .CK(clock), .Q(
        decode_regfile_fpregs_22__10_) );
  DFF_X2 decode_regfile_fpregs_reg_22__11_ ( .D(n7943), .CK(clock), .Q(
        decode_regfile_fpregs_22__11_) );
  DFF_X2 decode_regfile_fpregs_reg_22__12_ ( .D(n7942), .CK(clock), .Q(
        decode_regfile_fpregs_22__12_) );
  DFF_X2 decode_regfile_fpregs_reg_22__13_ ( .D(n7941), .CK(clock), .Q(
        decode_regfile_fpregs_22__13_) );
  DFF_X2 decode_regfile_fpregs_reg_22__14_ ( .D(n7940), .CK(clock), .Q(
        decode_regfile_fpregs_22__14_) );
  DFF_X2 decode_regfile_fpregs_reg_22__15_ ( .D(n7939), .CK(clock), .Q(
        decode_regfile_fpregs_22__15_) );
  DFF_X2 decode_regfile_fpregs_reg_22__16_ ( .D(n7938), .CK(clock), .Q(
        decode_regfile_fpregs_22__16_) );
  DFF_X2 decode_regfile_fpregs_reg_22__17_ ( .D(n7937), .CK(clock), .Q(
        decode_regfile_fpregs_22__17_) );
  DFF_X2 decode_regfile_fpregs_reg_22__18_ ( .D(n7936), .CK(clock), .Q(
        decode_regfile_fpregs_22__18_) );
  DFF_X2 decode_regfile_fpregs_reg_22__19_ ( .D(n7935), .CK(clock), .Q(
        decode_regfile_fpregs_22__19_) );
  DFF_X2 decode_regfile_fpregs_reg_22__20_ ( .D(n7934), .CK(clock), .Q(
        decode_regfile_fpregs_22__20_) );
  DFF_X2 decode_regfile_fpregs_reg_22__21_ ( .D(n7933), .CK(clock), .Q(
        decode_regfile_fpregs_22__21_) );
  DFF_X2 decode_regfile_fpregs_reg_22__22_ ( .D(n7932), .CK(clock), .Q(
        decode_regfile_fpregs_22__22_) );
  DFF_X2 decode_regfile_fpregs_reg_22__23_ ( .D(n7931), .CK(clock), .Q(
        decode_regfile_fpregs_22__23_) );
  DFF_X2 decode_regfile_fpregs_reg_22__24_ ( .D(n7930), .CK(clock), .Q(
        decode_regfile_fpregs_22__24_) );
  DFF_X2 decode_regfile_fpregs_reg_22__25_ ( .D(n7929), .CK(clock), .Q(
        decode_regfile_fpregs_22__25_) );
  DFF_X2 decode_regfile_fpregs_reg_22__26_ ( .D(n7928), .CK(clock), .Q(
        decode_regfile_fpregs_22__26_) );
  DFF_X2 decode_regfile_fpregs_reg_22__27_ ( .D(n7927), .CK(clock), .Q(
        decode_regfile_fpregs_22__27_) );
  DFF_X2 decode_regfile_fpregs_reg_22__28_ ( .D(n7926), .CK(clock), .Q(
        decode_regfile_fpregs_22__28_) );
  DFF_X2 decode_regfile_fpregs_reg_22__29_ ( .D(n7925), .CK(clock), .Q(
        decode_regfile_fpregs_22__29_) );
  DFF_X2 decode_regfile_fpregs_reg_22__30_ ( .D(n7924), .CK(clock), .Q(
        decode_regfile_fpregs_22__30_) );
  DFF_X2 decode_regfile_fpregs_reg_22__31_ ( .D(n7923), .CK(clock), .Q(
        decode_regfile_fpregs_22__31_) );
  DFF_X2 decode_regfile_fpregs_reg_21__0_ ( .D(n7922), .CK(clock), .Q(
        decode_regfile_fpregs_21__0_) );
  DFF_X2 decode_regfile_fpregs_reg_21__1_ ( .D(n7921), .CK(clock), .Q(
        decode_regfile_fpregs_21__1_) );
  DFF_X2 decode_regfile_fpregs_reg_21__2_ ( .D(n7920), .CK(clock), .Q(
        decode_regfile_fpregs_21__2_) );
  DFF_X2 decode_regfile_fpregs_reg_21__3_ ( .D(n7919), .CK(clock), .Q(
        decode_regfile_fpregs_21__3_) );
  DFF_X2 decode_regfile_fpregs_reg_21__4_ ( .D(n7918), .CK(clock), .Q(
        decode_regfile_fpregs_21__4_) );
  DFF_X2 decode_regfile_fpregs_reg_21__5_ ( .D(n7917), .CK(clock), .Q(
        decode_regfile_fpregs_21__5_) );
  DFF_X2 decode_regfile_fpregs_reg_21__6_ ( .D(n7916), .CK(clock), .Q(
        decode_regfile_fpregs_21__6_) );
  DFF_X2 decode_regfile_fpregs_reg_21__7_ ( .D(n7915), .CK(clock), .Q(
        decode_regfile_fpregs_21__7_) );
  DFF_X2 decode_regfile_fpregs_reg_21__8_ ( .D(n7914), .CK(clock), .Q(
        decode_regfile_fpregs_21__8_) );
  DFF_X2 decode_regfile_fpregs_reg_21__9_ ( .D(n7913), .CK(clock), .Q(
        decode_regfile_fpregs_21__9_) );
  DFF_X2 decode_regfile_fpregs_reg_21__10_ ( .D(n7912), .CK(clock), .Q(
        decode_regfile_fpregs_21__10_) );
  DFF_X2 decode_regfile_fpregs_reg_21__11_ ( .D(n7911), .CK(clock), .Q(
        decode_regfile_fpregs_21__11_) );
  DFF_X2 decode_regfile_fpregs_reg_21__12_ ( .D(n7910), .CK(clock), .Q(
        decode_regfile_fpregs_21__12_) );
  DFF_X2 decode_regfile_fpregs_reg_21__13_ ( .D(n7909), .CK(clock), .Q(
        decode_regfile_fpregs_21__13_) );
  DFF_X2 decode_regfile_fpregs_reg_21__14_ ( .D(n7908), .CK(clock), .Q(
        decode_regfile_fpregs_21__14_) );
  DFF_X2 decode_regfile_fpregs_reg_21__15_ ( .D(n7907), .CK(clock), .Q(
        decode_regfile_fpregs_21__15_) );
  DFF_X2 decode_regfile_fpregs_reg_21__16_ ( .D(n7906), .CK(clock), .Q(
        decode_regfile_fpregs_21__16_) );
  DFF_X2 decode_regfile_fpregs_reg_21__17_ ( .D(n7905), .CK(clock), .Q(
        decode_regfile_fpregs_21__17_) );
  DFF_X2 decode_regfile_fpregs_reg_21__18_ ( .D(n7904), .CK(clock), .Q(
        decode_regfile_fpregs_21__18_) );
  DFF_X2 decode_regfile_fpregs_reg_21__19_ ( .D(n7903), .CK(clock), .Q(
        decode_regfile_fpregs_21__19_) );
  DFF_X2 decode_regfile_fpregs_reg_21__20_ ( .D(n7902), .CK(clock), .Q(
        decode_regfile_fpregs_21__20_) );
  DFF_X2 decode_regfile_fpregs_reg_21__21_ ( .D(n7901), .CK(clock), .Q(
        decode_regfile_fpregs_21__21_) );
  DFF_X2 decode_regfile_fpregs_reg_21__22_ ( .D(n7900), .CK(clock), .Q(
        decode_regfile_fpregs_21__22_) );
  DFF_X2 decode_regfile_fpregs_reg_21__23_ ( .D(n7899), .CK(clock), .Q(
        decode_regfile_fpregs_21__23_) );
  DFF_X2 decode_regfile_fpregs_reg_21__24_ ( .D(n7898), .CK(clock), .Q(
        decode_regfile_fpregs_21__24_) );
  DFF_X2 decode_regfile_fpregs_reg_21__25_ ( .D(n7897), .CK(clock), .Q(
        decode_regfile_fpregs_21__25_) );
  DFF_X2 decode_regfile_fpregs_reg_21__26_ ( .D(n7896), .CK(clock), .Q(
        decode_regfile_fpregs_21__26_) );
  DFF_X2 decode_regfile_fpregs_reg_21__27_ ( .D(n7895), .CK(clock), .Q(
        decode_regfile_fpregs_21__27_) );
  DFF_X2 decode_regfile_fpregs_reg_21__28_ ( .D(n7894), .CK(clock), .Q(
        decode_regfile_fpregs_21__28_) );
  DFF_X2 decode_regfile_fpregs_reg_21__29_ ( .D(n7893), .CK(clock), .Q(
        decode_regfile_fpregs_21__29_) );
  DFF_X2 decode_regfile_fpregs_reg_21__30_ ( .D(n7892), .CK(clock), .Q(
        decode_regfile_fpregs_21__30_) );
  DFF_X2 decode_regfile_fpregs_reg_21__31_ ( .D(n7891), .CK(clock), .Q(
        decode_regfile_fpregs_21__31_) );
  DFF_X2 decode_regfile_fpregs_reg_20__0_ ( .D(n7890), .CK(clock), .Q(
        decode_regfile_fpregs_20__0_) );
  DFF_X2 decode_regfile_fpregs_reg_20__1_ ( .D(n7889), .CK(clock), .Q(
        decode_regfile_fpregs_20__1_) );
  DFF_X2 decode_regfile_fpregs_reg_20__2_ ( .D(n7888), .CK(clock), .Q(
        decode_regfile_fpregs_20__2_) );
  DFF_X2 decode_regfile_fpregs_reg_20__3_ ( .D(n7887), .CK(clock), .Q(
        decode_regfile_fpregs_20__3_) );
  DFF_X2 decode_regfile_fpregs_reg_20__4_ ( .D(n7886), .CK(clock), .Q(
        decode_regfile_fpregs_20__4_) );
  DFF_X2 decode_regfile_fpregs_reg_20__5_ ( .D(n7885), .CK(clock), .Q(
        decode_regfile_fpregs_20__5_) );
  DFF_X2 decode_regfile_fpregs_reg_20__6_ ( .D(n7884), .CK(clock), .Q(
        decode_regfile_fpregs_20__6_) );
  DFF_X2 decode_regfile_fpregs_reg_20__7_ ( .D(n7883), .CK(clock), .Q(
        decode_regfile_fpregs_20__7_) );
  DFF_X2 decode_regfile_fpregs_reg_20__8_ ( .D(n7882), .CK(clock), .Q(
        decode_regfile_fpregs_20__8_) );
  DFF_X2 decode_regfile_fpregs_reg_20__9_ ( .D(n7881), .CK(clock), .Q(
        decode_regfile_fpregs_20__9_) );
  DFF_X2 decode_regfile_fpregs_reg_20__10_ ( .D(n7880), .CK(clock), .Q(
        decode_regfile_fpregs_20__10_) );
  DFF_X2 decode_regfile_fpregs_reg_20__11_ ( .D(n7879), .CK(clock), .Q(
        decode_regfile_fpregs_20__11_) );
  DFF_X2 decode_regfile_fpregs_reg_20__12_ ( .D(n7878), .CK(clock), .Q(
        decode_regfile_fpregs_20__12_) );
  DFF_X2 decode_regfile_fpregs_reg_20__13_ ( .D(n7877), .CK(clock), .Q(
        decode_regfile_fpregs_20__13_) );
  DFF_X2 decode_regfile_fpregs_reg_20__14_ ( .D(n7876), .CK(clock), .Q(
        decode_regfile_fpregs_20__14_) );
  DFF_X2 decode_regfile_fpregs_reg_20__15_ ( .D(n7875), .CK(clock), .Q(
        decode_regfile_fpregs_20__15_) );
  DFF_X2 decode_regfile_fpregs_reg_20__16_ ( .D(n7874), .CK(clock), .Q(
        decode_regfile_fpregs_20__16_) );
  DFF_X2 decode_regfile_fpregs_reg_20__17_ ( .D(n7873), .CK(clock), .Q(
        decode_regfile_fpregs_20__17_) );
  DFF_X2 decode_regfile_fpregs_reg_20__18_ ( .D(n7872), .CK(clock), .Q(
        decode_regfile_fpregs_20__18_) );
  DFF_X2 decode_regfile_fpregs_reg_20__19_ ( .D(n7871), .CK(clock), .Q(
        decode_regfile_fpregs_20__19_) );
  DFF_X2 decode_regfile_fpregs_reg_20__20_ ( .D(n7870), .CK(clock), .Q(
        decode_regfile_fpregs_20__20_) );
  DFF_X2 decode_regfile_fpregs_reg_20__21_ ( .D(n7869), .CK(clock), .Q(
        decode_regfile_fpregs_20__21_) );
  DFF_X2 decode_regfile_fpregs_reg_20__22_ ( .D(n7868), .CK(clock), .Q(
        decode_regfile_fpregs_20__22_) );
  DFF_X2 decode_regfile_fpregs_reg_20__23_ ( .D(n7867), .CK(clock), .Q(
        decode_regfile_fpregs_20__23_) );
  DFF_X2 decode_regfile_fpregs_reg_20__24_ ( .D(n7866), .CK(clock), .Q(
        decode_regfile_fpregs_20__24_) );
  DFF_X2 decode_regfile_fpregs_reg_20__25_ ( .D(n7865), .CK(clock), .Q(
        decode_regfile_fpregs_20__25_) );
  DFF_X2 decode_regfile_fpregs_reg_20__26_ ( .D(n7864), .CK(clock), .Q(
        decode_regfile_fpregs_20__26_) );
  DFF_X2 decode_regfile_fpregs_reg_20__27_ ( .D(n7863), .CK(clock), .Q(
        decode_regfile_fpregs_20__27_) );
  DFF_X2 decode_regfile_fpregs_reg_20__28_ ( .D(n7862), .CK(clock), .Q(
        decode_regfile_fpregs_20__28_) );
  DFF_X2 decode_regfile_fpregs_reg_20__29_ ( .D(n7861), .CK(clock), .Q(
        decode_regfile_fpregs_20__29_) );
  DFF_X2 decode_regfile_fpregs_reg_20__30_ ( .D(n7860), .CK(clock), .Q(
        decode_regfile_fpregs_20__30_) );
  DFF_X2 decode_regfile_fpregs_reg_20__31_ ( .D(n7859), .CK(clock), .Q(
        decode_regfile_fpregs_20__31_) );
  DFF_X2 decode_regfile_fpregs_reg_19__0_ ( .D(n7858), .CK(clock), .Q(
        decode_regfile_fpregs_19__0_) );
  DFF_X2 decode_regfile_fpregs_reg_19__1_ ( .D(n7857), .CK(clock), .Q(
        decode_regfile_fpregs_19__1_) );
  DFF_X2 decode_regfile_fpregs_reg_19__2_ ( .D(n7856), .CK(clock), .Q(
        decode_regfile_fpregs_19__2_) );
  DFF_X2 decode_regfile_fpregs_reg_19__3_ ( .D(n7855), .CK(clock), .Q(
        decode_regfile_fpregs_19__3_) );
  DFF_X2 decode_regfile_fpregs_reg_19__4_ ( .D(n7854), .CK(clock), .Q(
        decode_regfile_fpregs_19__4_) );
  DFF_X2 decode_regfile_fpregs_reg_19__5_ ( .D(n7853), .CK(clock), .Q(
        decode_regfile_fpregs_19__5_) );
  DFF_X2 decode_regfile_fpregs_reg_19__6_ ( .D(n7852), .CK(clock), .Q(
        decode_regfile_fpregs_19__6_) );
  DFF_X2 decode_regfile_fpregs_reg_19__7_ ( .D(n7851), .CK(clock), .Q(
        decode_regfile_fpregs_19__7_) );
  DFF_X2 decode_regfile_fpregs_reg_19__8_ ( .D(n7850), .CK(clock), .Q(
        decode_regfile_fpregs_19__8_) );
  DFF_X2 decode_regfile_fpregs_reg_19__9_ ( .D(n7849), .CK(clock), .Q(
        decode_regfile_fpregs_19__9_) );
  DFF_X2 decode_regfile_fpregs_reg_19__10_ ( .D(n7848), .CK(clock), .Q(
        decode_regfile_fpregs_19__10_) );
  DFF_X2 decode_regfile_fpregs_reg_19__11_ ( .D(n7847), .CK(clock), .Q(
        decode_regfile_fpregs_19__11_) );
  DFF_X2 decode_regfile_fpregs_reg_19__12_ ( .D(n7846), .CK(clock), .Q(
        decode_regfile_fpregs_19__12_) );
  DFF_X2 decode_regfile_fpregs_reg_19__13_ ( .D(n7845), .CK(clock), .Q(
        decode_regfile_fpregs_19__13_) );
  DFF_X2 decode_regfile_fpregs_reg_19__14_ ( .D(n7844), .CK(clock), .Q(
        decode_regfile_fpregs_19__14_) );
  DFF_X2 decode_regfile_fpregs_reg_19__15_ ( .D(n7843), .CK(clock), .Q(
        decode_regfile_fpregs_19__15_) );
  DFF_X2 decode_regfile_fpregs_reg_19__16_ ( .D(n7842), .CK(clock), .Q(
        decode_regfile_fpregs_19__16_) );
  DFF_X2 decode_regfile_fpregs_reg_19__17_ ( .D(n7841), .CK(clock), .Q(
        decode_regfile_fpregs_19__17_) );
  DFF_X2 decode_regfile_fpregs_reg_19__18_ ( .D(n7840), .CK(clock), .Q(
        decode_regfile_fpregs_19__18_) );
  DFF_X2 decode_regfile_fpregs_reg_19__19_ ( .D(n7839), .CK(clock), .Q(
        decode_regfile_fpregs_19__19_) );
  DFF_X2 decode_regfile_fpregs_reg_19__20_ ( .D(n7838), .CK(clock), .Q(
        decode_regfile_fpregs_19__20_) );
  DFF_X2 decode_regfile_fpregs_reg_19__21_ ( .D(n7837), .CK(clock), .Q(
        decode_regfile_fpregs_19__21_) );
  DFF_X2 decode_regfile_fpregs_reg_19__22_ ( .D(n7836), .CK(clock), .Q(
        decode_regfile_fpregs_19__22_) );
  DFF_X2 decode_regfile_fpregs_reg_19__23_ ( .D(n7835), .CK(clock), .Q(
        decode_regfile_fpregs_19__23_) );
  DFF_X2 decode_regfile_fpregs_reg_19__24_ ( .D(n7834), .CK(clock), .Q(
        decode_regfile_fpregs_19__24_) );
  DFF_X2 decode_regfile_fpregs_reg_19__25_ ( .D(n7833), .CK(clock), .Q(
        decode_regfile_fpregs_19__25_) );
  DFF_X2 decode_regfile_fpregs_reg_19__26_ ( .D(n7832), .CK(clock), .Q(
        decode_regfile_fpregs_19__26_) );
  DFF_X2 decode_regfile_fpregs_reg_19__27_ ( .D(n7831), .CK(clock), .Q(
        decode_regfile_fpregs_19__27_) );
  DFF_X2 decode_regfile_fpregs_reg_19__28_ ( .D(n7830), .CK(clock), .Q(
        decode_regfile_fpregs_19__28_) );
  DFF_X2 decode_regfile_fpregs_reg_19__29_ ( .D(n7829), .CK(clock), .Q(
        decode_regfile_fpregs_19__29_) );
  DFF_X2 decode_regfile_fpregs_reg_19__30_ ( .D(n7828), .CK(clock), .Q(
        decode_regfile_fpregs_19__30_) );
  DFF_X2 decode_regfile_fpregs_reg_19__31_ ( .D(n7827), .CK(clock), .Q(
        decode_regfile_fpregs_19__31_) );
  DFF_X2 decode_regfile_fpregs_reg_18__0_ ( .D(n7826), .CK(clock), .Q(
        decode_regfile_fpregs_18__0_) );
  DFF_X2 decode_regfile_fpregs_reg_18__1_ ( .D(n7825), .CK(clock), .Q(
        decode_regfile_fpregs_18__1_) );
  DFF_X2 decode_regfile_fpregs_reg_18__2_ ( .D(n7824), .CK(clock), .Q(
        decode_regfile_fpregs_18__2_) );
  DFF_X2 decode_regfile_fpregs_reg_18__3_ ( .D(n7823), .CK(clock), .Q(
        decode_regfile_fpregs_18__3_) );
  DFF_X2 decode_regfile_fpregs_reg_18__4_ ( .D(n7822), .CK(clock), .Q(
        decode_regfile_fpregs_18__4_) );
  DFF_X2 decode_regfile_fpregs_reg_18__5_ ( .D(n7821), .CK(clock), .Q(
        decode_regfile_fpregs_18__5_) );
  DFF_X2 decode_regfile_fpregs_reg_18__6_ ( .D(n7820), .CK(clock), .Q(
        decode_regfile_fpregs_18__6_) );
  DFF_X2 decode_regfile_fpregs_reg_18__7_ ( .D(n7819), .CK(clock), .Q(
        decode_regfile_fpregs_18__7_) );
  DFF_X2 decode_regfile_fpregs_reg_18__8_ ( .D(n7818), .CK(clock), .Q(
        decode_regfile_fpregs_18__8_) );
  DFF_X2 decode_regfile_fpregs_reg_18__9_ ( .D(n7817), .CK(clock), .Q(
        decode_regfile_fpregs_18__9_) );
  DFF_X2 decode_regfile_fpregs_reg_18__10_ ( .D(n7816), .CK(clock), .Q(
        decode_regfile_fpregs_18__10_) );
  DFF_X2 decode_regfile_fpregs_reg_18__11_ ( .D(n7815), .CK(clock), .Q(
        decode_regfile_fpregs_18__11_) );
  DFF_X2 decode_regfile_fpregs_reg_18__12_ ( .D(n7814), .CK(clock), .Q(
        decode_regfile_fpregs_18__12_) );
  DFF_X2 decode_regfile_fpregs_reg_18__13_ ( .D(n7813), .CK(clock), .Q(
        decode_regfile_fpregs_18__13_) );
  DFF_X2 decode_regfile_fpregs_reg_18__14_ ( .D(n7812), .CK(clock), .Q(
        decode_regfile_fpregs_18__14_) );
  DFF_X2 decode_regfile_fpregs_reg_18__15_ ( .D(n7811), .CK(clock), .Q(
        decode_regfile_fpregs_18__15_) );
  DFF_X2 decode_regfile_fpregs_reg_18__16_ ( .D(n7810), .CK(clock), .Q(
        decode_regfile_fpregs_18__16_) );
  DFF_X2 decode_regfile_fpregs_reg_18__17_ ( .D(n7809), .CK(clock), .Q(
        decode_regfile_fpregs_18__17_) );
  DFF_X2 decode_regfile_fpregs_reg_18__18_ ( .D(n7808), .CK(clock), .Q(
        decode_regfile_fpregs_18__18_) );
  DFF_X2 decode_regfile_fpregs_reg_18__19_ ( .D(n7807), .CK(clock), .Q(
        decode_regfile_fpregs_18__19_) );
  DFF_X2 decode_regfile_fpregs_reg_18__20_ ( .D(n7806), .CK(clock), .Q(
        decode_regfile_fpregs_18__20_) );
  DFF_X2 decode_regfile_fpregs_reg_18__21_ ( .D(n7805), .CK(clock), .Q(
        decode_regfile_fpregs_18__21_) );
  DFF_X2 decode_regfile_fpregs_reg_18__22_ ( .D(n7804), .CK(clock), .Q(
        decode_regfile_fpregs_18__22_) );
  DFF_X2 decode_regfile_fpregs_reg_18__23_ ( .D(n7803), .CK(clock), .Q(
        decode_regfile_fpregs_18__23_) );
  DFF_X2 decode_regfile_fpregs_reg_18__24_ ( .D(n7802), .CK(clock), .Q(
        decode_regfile_fpregs_18__24_) );
  DFF_X2 decode_regfile_fpregs_reg_18__25_ ( .D(n7801), .CK(clock), .Q(
        decode_regfile_fpregs_18__25_) );
  DFF_X2 decode_regfile_fpregs_reg_18__26_ ( .D(n7800), .CK(clock), .Q(
        decode_regfile_fpregs_18__26_) );
  DFF_X2 decode_regfile_fpregs_reg_18__27_ ( .D(n7799), .CK(clock), .Q(
        decode_regfile_fpregs_18__27_) );
  DFF_X2 decode_regfile_fpregs_reg_18__28_ ( .D(n7798), .CK(clock), .Q(
        decode_regfile_fpregs_18__28_) );
  DFF_X2 decode_regfile_fpregs_reg_18__29_ ( .D(n7797), .CK(clock), .Q(
        decode_regfile_fpregs_18__29_) );
  DFF_X2 decode_regfile_fpregs_reg_18__30_ ( .D(n7796), .CK(clock), .Q(
        decode_regfile_fpregs_18__30_) );
  DFF_X2 decode_regfile_fpregs_reg_18__31_ ( .D(n7795), .CK(clock), .Q(
        decode_regfile_fpregs_18__31_) );
  DFF_X2 decode_regfile_fpregs_reg_17__0_ ( .D(n7794), .CK(clock), .Q(
        decode_regfile_fpregs_17__0_) );
  DFF_X2 decode_regfile_fpregs_reg_17__1_ ( .D(n7793), .CK(clock), .Q(
        decode_regfile_fpregs_17__1_) );
  DFF_X2 decode_regfile_fpregs_reg_17__2_ ( .D(n7792), .CK(clock), .Q(
        decode_regfile_fpregs_17__2_) );
  DFF_X2 decode_regfile_fpregs_reg_17__3_ ( .D(n7791), .CK(clock), .Q(
        decode_regfile_fpregs_17__3_) );
  DFF_X2 decode_regfile_fpregs_reg_17__4_ ( .D(n7790), .CK(clock), .Q(
        decode_regfile_fpregs_17__4_) );
  DFF_X2 decode_regfile_fpregs_reg_17__5_ ( .D(n7789), .CK(clock), .Q(
        decode_regfile_fpregs_17__5_) );
  DFF_X2 decode_regfile_fpregs_reg_17__6_ ( .D(n7788), .CK(clock), .Q(
        decode_regfile_fpregs_17__6_) );
  DFF_X2 decode_regfile_fpregs_reg_17__7_ ( .D(n7787), .CK(clock), .Q(
        decode_regfile_fpregs_17__7_) );
  DFF_X2 decode_regfile_fpregs_reg_17__8_ ( .D(n7786), .CK(clock), .Q(
        decode_regfile_fpregs_17__8_) );
  DFF_X2 decode_regfile_fpregs_reg_17__9_ ( .D(n7785), .CK(clock), .Q(
        decode_regfile_fpregs_17__9_) );
  DFF_X2 decode_regfile_fpregs_reg_17__10_ ( .D(n7784), .CK(clock), .Q(
        decode_regfile_fpregs_17__10_) );
  DFF_X2 decode_regfile_fpregs_reg_17__11_ ( .D(n7783), .CK(clock), .Q(
        decode_regfile_fpregs_17__11_) );
  DFF_X2 decode_regfile_fpregs_reg_17__12_ ( .D(n7782), .CK(clock), .Q(
        decode_regfile_fpregs_17__12_) );
  DFF_X2 decode_regfile_fpregs_reg_17__13_ ( .D(n7781), .CK(clock), .Q(
        decode_regfile_fpregs_17__13_) );
  DFF_X2 decode_regfile_fpregs_reg_17__14_ ( .D(n7780), .CK(clock), .Q(
        decode_regfile_fpregs_17__14_) );
  DFF_X2 decode_regfile_fpregs_reg_17__15_ ( .D(n7779), .CK(clock), .Q(
        decode_regfile_fpregs_17__15_) );
  DFF_X2 decode_regfile_fpregs_reg_17__16_ ( .D(n7778), .CK(clock), .Q(
        decode_regfile_fpregs_17__16_) );
  DFF_X2 decode_regfile_fpregs_reg_17__17_ ( .D(n7777), .CK(clock), .Q(
        decode_regfile_fpregs_17__17_) );
  DFF_X2 decode_regfile_fpregs_reg_17__18_ ( .D(n7776), .CK(clock), .Q(
        decode_regfile_fpregs_17__18_) );
  DFF_X2 decode_regfile_fpregs_reg_17__19_ ( .D(n7775), .CK(clock), .Q(
        decode_regfile_fpregs_17__19_) );
  DFF_X2 decode_regfile_fpregs_reg_17__20_ ( .D(n7774), .CK(clock), .Q(
        decode_regfile_fpregs_17__20_) );
  DFF_X2 decode_regfile_fpregs_reg_17__21_ ( .D(n7773), .CK(clock), .Q(
        decode_regfile_fpregs_17__21_) );
  DFF_X2 decode_regfile_fpregs_reg_17__22_ ( .D(n7772), .CK(clock), .Q(
        decode_regfile_fpregs_17__22_) );
  DFF_X2 decode_regfile_fpregs_reg_17__23_ ( .D(n7771), .CK(clock), .Q(
        decode_regfile_fpregs_17__23_) );
  DFF_X2 decode_regfile_fpregs_reg_17__24_ ( .D(n7770), .CK(clock), .Q(
        decode_regfile_fpregs_17__24_) );
  DFF_X2 decode_regfile_fpregs_reg_17__25_ ( .D(n7769), .CK(clock), .Q(
        decode_regfile_fpregs_17__25_) );
  DFF_X2 decode_regfile_fpregs_reg_17__26_ ( .D(n7768), .CK(clock), .Q(
        decode_regfile_fpregs_17__26_) );
  DFF_X2 decode_regfile_fpregs_reg_17__27_ ( .D(n7767), .CK(clock), .Q(
        decode_regfile_fpregs_17__27_) );
  DFF_X2 decode_regfile_fpregs_reg_17__28_ ( .D(n7766), .CK(clock), .Q(
        decode_regfile_fpregs_17__28_) );
  DFF_X2 decode_regfile_fpregs_reg_17__29_ ( .D(n7765), .CK(clock), .Q(
        decode_regfile_fpregs_17__29_) );
  DFF_X2 decode_regfile_fpregs_reg_17__30_ ( .D(n7764), .CK(clock), .Q(
        decode_regfile_fpregs_17__30_) );
  DFF_X2 decode_regfile_fpregs_reg_17__31_ ( .D(n7763), .CK(clock), .Q(
        decode_regfile_fpregs_17__31_) );
  DFF_X2 decode_regfile_fpregs_reg_16__0_ ( .D(n7762), .CK(clock), .Q(
        decode_regfile_fpregs_16__0_) );
  DFF_X2 decode_regfile_fpregs_reg_16__1_ ( .D(n7761), .CK(clock), .Q(
        decode_regfile_fpregs_16__1_) );
  DFF_X2 decode_regfile_fpregs_reg_16__2_ ( .D(n7760), .CK(clock), .Q(
        decode_regfile_fpregs_16__2_) );
  DFF_X2 decode_regfile_fpregs_reg_16__3_ ( .D(n7759), .CK(clock), .Q(
        decode_regfile_fpregs_16__3_) );
  DFF_X2 decode_regfile_fpregs_reg_16__4_ ( .D(n7758), .CK(clock), .Q(
        decode_regfile_fpregs_16__4_) );
  DFF_X2 decode_regfile_fpregs_reg_16__5_ ( .D(n7757), .CK(clock), .Q(
        decode_regfile_fpregs_16__5_) );
  DFF_X2 decode_regfile_fpregs_reg_16__6_ ( .D(n7756), .CK(clock), .Q(
        decode_regfile_fpregs_16__6_) );
  DFF_X2 decode_regfile_fpregs_reg_16__7_ ( .D(n7755), .CK(clock), .Q(
        decode_regfile_fpregs_16__7_) );
  DFF_X2 decode_regfile_fpregs_reg_16__8_ ( .D(n7754), .CK(clock), .Q(
        decode_regfile_fpregs_16__8_) );
  DFF_X2 decode_regfile_fpregs_reg_16__9_ ( .D(n7753), .CK(clock), .Q(
        decode_regfile_fpregs_16__9_) );
  DFF_X2 decode_regfile_fpregs_reg_16__10_ ( .D(n7752), .CK(clock), .Q(
        decode_regfile_fpregs_16__10_) );
  DFF_X2 decode_regfile_fpregs_reg_16__11_ ( .D(n7751), .CK(clock), .Q(
        decode_regfile_fpregs_16__11_) );
  DFF_X2 decode_regfile_fpregs_reg_16__12_ ( .D(n7750), .CK(clock), .Q(
        decode_regfile_fpregs_16__12_) );
  DFF_X2 decode_regfile_fpregs_reg_16__13_ ( .D(n7749), .CK(clock), .Q(
        decode_regfile_fpregs_16__13_) );
  DFF_X2 decode_regfile_fpregs_reg_16__14_ ( .D(n7748), .CK(clock), .Q(
        decode_regfile_fpregs_16__14_) );
  DFF_X2 decode_regfile_fpregs_reg_16__15_ ( .D(n7747), .CK(clock), .Q(
        decode_regfile_fpregs_16__15_) );
  DFF_X2 decode_regfile_fpregs_reg_16__16_ ( .D(n7746), .CK(clock), .Q(
        decode_regfile_fpregs_16__16_) );
  DFF_X2 decode_regfile_fpregs_reg_16__17_ ( .D(n7745), .CK(clock), .Q(
        decode_regfile_fpregs_16__17_) );
  DFF_X2 decode_regfile_fpregs_reg_16__18_ ( .D(n7744), .CK(clock), .Q(
        decode_regfile_fpregs_16__18_) );
  DFF_X2 decode_regfile_fpregs_reg_16__19_ ( .D(n7743), .CK(clock), .Q(
        decode_regfile_fpregs_16__19_) );
  DFF_X2 decode_regfile_fpregs_reg_16__20_ ( .D(n7742), .CK(clock), .Q(
        decode_regfile_fpregs_16__20_) );
  DFF_X2 decode_regfile_fpregs_reg_16__21_ ( .D(n7741), .CK(clock), .Q(
        decode_regfile_fpregs_16__21_) );
  DFF_X2 decode_regfile_fpregs_reg_16__22_ ( .D(n7740), .CK(clock), .Q(
        decode_regfile_fpregs_16__22_) );
  DFF_X2 decode_regfile_fpregs_reg_16__23_ ( .D(n7739), .CK(clock), .Q(
        decode_regfile_fpregs_16__23_) );
  DFF_X2 decode_regfile_fpregs_reg_16__24_ ( .D(n7738), .CK(clock), .Q(
        decode_regfile_fpregs_16__24_) );
  DFF_X2 decode_regfile_fpregs_reg_16__25_ ( .D(n7737), .CK(clock), .Q(
        decode_regfile_fpregs_16__25_) );
  DFF_X2 decode_regfile_fpregs_reg_16__26_ ( .D(n7736), .CK(clock), .Q(
        decode_regfile_fpregs_16__26_) );
  DFF_X2 decode_regfile_fpregs_reg_16__27_ ( .D(n7735), .CK(clock), .Q(
        decode_regfile_fpregs_16__27_) );
  DFF_X2 decode_regfile_fpregs_reg_16__28_ ( .D(n7734), .CK(clock), .Q(
        decode_regfile_fpregs_16__28_) );
  DFF_X2 decode_regfile_fpregs_reg_16__29_ ( .D(n7733), .CK(clock), .Q(
        decode_regfile_fpregs_16__29_) );
  DFF_X2 decode_regfile_fpregs_reg_16__30_ ( .D(n7732), .CK(clock), .Q(
        decode_regfile_fpregs_16__30_) );
  DFF_X2 decode_regfile_fpregs_reg_16__31_ ( .D(n7731), .CK(clock), .Q(
        decode_regfile_fpregs_16__31_) );
  DFF_X2 decode_regfile_fpregs_reg_15__0_ ( .D(n7730), .CK(clock), .Q(
        decode_regfile_fpregs_15__0_) );
  DFF_X2 decode_regfile_fpregs_reg_15__1_ ( .D(n7729), .CK(clock), .Q(
        decode_regfile_fpregs_15__1_) );
  DFF_X2 decode_regfile_fpregs_reg_15__2_ ( .D(n7728), .CK(clock), .Q(
        decode_regfile_fpregs_15__2_) );
  DFF_X2 decode_regfile_fpregs_reg_15__3_ ( .D(n7727), .CK(clock), .Q(
        decode_regfile_fpregs_15__3_) );
  DFF_X2 decode_regfile_fpregs_reg_15__4_ ( .D(n7726), .CK(clock), .Q(
        decode_regfile_fpregs_15__4_) );
  DFF_X2 decode_regfile_fpregs_reg_15__5_ ( .D(n7725), .CK(clock), .Q(
        decode_regfile_fpregs_15__5_) );
  DFF_X2 decode_regfile_fpregs_reg_15__6_ ( .D(n7724), .CK(clock), .Q(
        decode_regfile_fpregs_15__6_) );
  DFF_X2 decode_regfile_fpregs_reg_15__7_ ( .D(n7723), .CK(clock), .Q(
        decode_regfile_fpregs_15__7_) );
  DFF_X2 decode_regfile_fpregs_reg_15__8_ ( .D(n7722), .CK(clock), .Q(
        decode_regfile_fpregs_15__8_) );
  DFF_X2 decode_regfile_fpregs_reg_15__9_ ( .D(n7721), .CK(clock), .Q(
        decode_regfile_fpregs_15__9_) );
  DFF_X2 decode_regfile_fpregs_reg_15__10_ ( .D(n7720), .CK(clock), .Q(
        decode_regfile_fpregs_15__10_) );
  DFF_X2 decode_regfile_fpregs_reg_15__11_ ( .D(n7719), .CK(clock), .Q(
        decode_regfile_fpregs_15__11_) );
  DFF_X2 decode_regfile_fpregs_reg_15__12_ ( .D(n7718), .CK(clock), .Q(
        decode_regfile_fpregs_15__12_) );
  DFF_X2 decode_regfile_fpregs_reg_15__13_ ( .D(n7717), .CK(clock), .Q(
        decode_regfile_fpregs_15__13_) );
  DFF_X2 decode_regfile_fpregs_reg_15__14_ ( .D(n7716), .CK(clock), .Q(
        decode_regfile_fpregs_15__14_) );
  DFF_X2 decode_regfile_fpregs_reg_15__15_ ( .D(n7715), .CK(clock), .Q(
        decode_regfile_fpregs_15__15_) );
  DFF_X2 decode_regfile_fpregs_reg_15__16_ ( .D(n7714), .CK(clock), .Q(
        decode_regfile_fpregs_15__16_) );
  DFF_X2 decode_regfile_fpregs_reg_15__17_ ( .D(n7713), .CK(clock), .Q(
        decode_regfile_fpregs_15__17_) );
  DFF_X2 decode_regfile_fpregs_reg_15__18_ ( .D(n7712), .CK(clock), .Q(
        decode_regfile_fpregs_15__18_) );
  DFF_X2 decode_regfile_fpregs_reg_15__19_ ( .D(n7711), .CK(clock), .Q(
        decode_regfile_fpregs_15__19_) );
  DFF_X2 decode_regfile_fpregs_reg_15__20_ ( .D(n7710), .CK(clock), .Q(
        decode_regfile_fpregs_15__20_) );
  DFF_X2 decode_regfile_fpregs_reg_15__21_ ( .D(n7709), .CK(clock), .Q(
        decode_regfile_fpregs_15__21_) );
  DFF_X2 decode_regfile_fpregs_reg_15__22_ ( .D(n7708), .CK(clock), .Q(
        decode_regfile_fpregs_15__22_) );
  DFF_X2 decode_regfile_fpregs_reg_15__23_ ( .D(n7707), .CK(clock), .Q(
        decode_regfile_fpregs_15__23_) );
  DFF_X2 decode_regfile_fpregs_reg_15__24_ ( .D(n7706), .CK(clock), .Q(
        decode_regfile_fpregs_15__24_) );
  DFF_X2 decode_regfile_fpregs_reg_15__25_ ( .D(n7705), .CK(clock), .Q(
        decode_regfile_fpregs_15__25_) );
  DFF_X2 decode_regfile_fpregs_reg_15__26_ ( .D(n7704), .CK(clock), .Q(
        decode_regfile_fpregs_15__26_) );
  DFF_X2 decode_regfile_fpregs_reg_15__27_ ( .D(n7703), .CK(clock), .Q(
        decode_regfile_fpregs_15__27_) );
  DFF_X2 decode_regfile_fpregs_reg_15__28_ ( .D(n7702), .CK(clock), .Q(
        decode_regfile_fpregs_15__28_) );
  DFF_X2 decode_regfile_fpregs_reg_15__29_ ( .D(n7701), .CK(clock), .Q(
        decode_regfile_fpregs_15__29_) );
  DFF_X2 decode_regfile_fpregs_reg_15__30_ ( .D(n7700), .CK(clock), .Q(
        decode_regfile_fpregs_15__30_) );
  DFF_X2 decode_regfile_fpregs_reg_15__31_ ( .D(n7699), .CK(clock), .Q(
        decode_regfile_fpregs_15__31_) );
  DFF_X2 decode_regfile_fpregs_reg_14__0_ ( .D(n7698), .CK(clock), .Q(
        decode_regfile_fpregs_14__0_) );
  DFF_X2 decode_regfile_fpregs_reg_14__1_ ( .D(n7697), .CK(clock), .Q(
        decode_regfile_fpregs_14__1_) );
  DFF_X2 decode_regfile_fpregs_reg_14__2_ ( .D(n7696), .CK(clock), .Q(
        decode_regfile_fpregs_14__2_) );
  DFF_X2 decode_regfile_fpregs_reg_14__3_ ( .D(n7695), .CK(clock), .Q(
        decode_regfile_fpregs_14__3_) );
  DFF_X2 decode_regfile_fpregs_reg_14__4_ ( .D(n7694), .CK(clock), .Q(
        decode_regfile_fpregs_14__4_) );
  DFF_X2 decode_regfile_fpregs_reg_14__5_ ( .D(n7693), .CK(clock), .Q(
        decode_regfile_fpregs_14__5_) );
  DFF_X2 decode_regfile_fpregs_reg_14__6_ ( .D(n7692), .CK(clock), .Q(
        decode_regfile_fpregs_14__6_) );
  DFF_X2 decode_regfile_fpregs_reg_14__7_ ( .D(n7691), .CK(clock), .Q(
        decode_regfile_fpregs_14__7_) );
  DFF_X2 decode_regfile_fpregs_reg_14__8_ ( .D(n7690), .CK(clock), .Q(
        decode_regfile_fpregs_14__8_) );
  DFF_X2 decode_regfile_fpregs_reg_14__9_ ( .D(n7689), .CK(clock), .Q(
        decode_regfile_fpregs_14__9_) );
  DFF_X2 decode_regfile_fpregs_reg_14__10_ ( .D(n7688), .CK(clock), .Q(
        decode_regfile_fpregs_14__10_) );
  DFF_X2 decode_regfile_fpregs_reg_14__11_ ( .D(n7687), .CK(clock), .Q(
        decode_regfile_fpregs_14__11_) );
  DFF_X2 decode_regfile_fpregs_reg_14__12_ ( .D(n7686), .CK(clock), .Q(
        decode_regfile_fpregs_14__12_) );
  DFF_X2 decode_regfile_fpregs_reg_14__13_ ( .D(n7685), .CK(clock), .Q(
        decode_regfile_fpregs_14__13_) );
  DFF_X2 decode_regfile_fpregs_reg_14__14_ ( .D(n7684), .CK(clock), .Q(
        decode_regfile_fpregs_14__14_) );
  DFF_X2 decode_regfile_fpregs_reg_14__15_ ( .D(n7683), .CK(clock), .Q(
        decode_regfile_fpregs_14__15_) );
  DFF_X2 decode_regfile_fpregs_reg_14__16_ ( .D(n7682), .CK(clock), .Q(
        decode_regfile_fpregs_14__16_) );
  DFF_X2 decode_regfile_fpregs_reg_14__17_ ( .D(n7681), .CK(clock), .Q(
        decode_regfile_fpregs_14__17_) );
  DFF_X2 decode_regfile_fpregs_reg_14__18_ ( .D(n7680), .CK(clock), .Q(
        decode_regfile_fpregs_14__18_) );
  DFF_X2 decode_regfile_fpregs_reg_14__19_ ( .D(n7679), .CK(clock), .Q(
        decode_regfile_fpregs_14__19_) );
  DFF_X2 decode_regfile_fpregs_reg_14__20_ ( .D(n7678), .CK(clock), .Q(
        decode_regfile_fpregs_14__20_) );
  DFF_X2 decode_regfile_fpregs_reg_14__21_ ( .D(n7677), .CK(clock), .Q(
        decode_regfile_fpregs_14__21_) );
  DFF_X2 decode_regfile_fpregs_reg_14__22_ ( .D(n7676), .CK(clock), .Q(
        decode_regfile_fpregs_14__22_) );
  DFF_X2 decode_regfile_fpregs_reg_14__23_ ( .D(n7675), .CK(clock), .Q(
        decode_regfile_fpregs_14__23_) );
  DFF_X2 decode_regfile_fpregs_reg_14__24_ ( .D(n7674), .CK(clock), .Q(
        decode_regfile_fpregs_14__24_) );
  DFF_X2 decode_regfile_fpregs_reg_14__25_ ( .D(n7673), .CK(clock), .Q(
        decode_regfile_fpregs_14__25_) );
  DFF_X2 decode_regfile_fpregs_reg_14__26_ ( .D(n7672), .CK(clock), .Q(
        decode_regfile_fpregs_14__26_) );
  DFF_X2 decode_regfile_fpregs_reg_14__27_ ( .D(n7671), .CK(clock), .Q(
        decode_regfile_fpregs_14__27_) );
  DFF_X2 decode_regfile_fpregs_reg_14__28_ ( .D(n7670), .CK(clock), .Q(
        decode_regfile_fpregs_14__28_) );
  DFF_X2 decode_regfile_fpregs_reg_14__29_ ( .D(n7669), .CK(clock), .Q(
        decode_regfile_fpregs_14__29_) );
  DFF_X2 decode_regfile_fpregs_reg_14__30_ ( .D(n7668), .CK(clock), .Q(
        decode_regfile_fpregs_14__30_) );
  DFF_X2 decode_regfile_fpregs_reg_14__31_ ( .D(n7667), .CK(clock), .Q(
        decode_regfile_fpregs_14__31_) );
  DFF_X2 decode_regfile_fpregs_reg_13__0_ ( .D(n7666), .CK(clock), .Q(
        decode_regfile_fpregs_13__0_) );
  DFF_X2 decode_regfile_fpregs_reg_13__1_ ( .D(n7665), .CK(clock), .Q(
        decode_regfile_fpregs_13__1_) );
  DFF_X2 decode_regfile_fpregs_reg_13__2_ ( .D(n7664), .CK(clock), .Q(
        decode_regfile_fpregs_13__2_) );
  DFF_X2 decode_regfile_fpregs_reg_13__3_ ( .D(n7663), .CK(clock), .Q(
        decode_regfile_fpregs_13__3_) );
  DFF_X2 decode_regfile_fpregs_reg_13__4_ ( .D(n7662), .CK(clock), .Q(
        decode_regfile_fpregs_13__4_) );
  DFF_X2 decode_regfile_fpregs_reg_13__5_ ( .D(n7661), .CK(clock), .Q(
        decode_regfile_fpregs_13__5_) );
  DFF_X2 decode_regfile_fpregs_reg_13__6_ ( .D(n7660), .CK(clock), .Q(
        decode_regfile_fpregs_13__6_) );
  DFF_X2 decode_regfile_fpregs_reg_13__7_ ( .D(n7659), .CK(clock), .Q(
        decode_regfile_fpregs_13__7_) );
  DFF_X2 decode_regfile_fpregs_reg_13__8_ ( .D(n7658), .CK(clock), .Q(
        decode_regfile_fpregs_13__8_) );
  DFF_X2 decode_regfile_fpregs_reg_13__9_ ( .D(n7657), .CK(clock), .Q(
        decode_regfile_fpregs_13__9_) );
  DFF_X2 decode_regfile_fpregs_reg_13__10_ ( .D(n7656), .CK(clock), .Q(
        decode_regfile_fpregs_13__10_) );
  DFF_X2 decode_regfile_fpregs_reg_13__11_ ( .D(n7655), .CK(clock), .Q(
        decode_regfile_fpregs_13__11_) );
  DFF_X2 decode_regfile_fpregs_reg_13__12_ ( .D(n7654), .CK(clock), .Q(
        decode_regfile_fpregs_13__12_) );
  DFF_X2 decode_regfile_fpregs_reg_13__13_ ( .D(n7653), .CK(clock), .Q(
        decode_regfile_fpregs_13__13_) );
  DFF_X2 decode_regfile_fpregs_reg_13__14_ ( .D(n7652), .CK(clock), .Q(
        decode_regfile_fpregs_13__14_) );
  DFF_X2 decode_regfile_fpregs_reg_13__15_ ( .D(n7651), .CK(clock), .Q(
        decode_regfile_fpregs_13__15_) );
  DFF_X2 decode_regfile_fpregs_reg_13__16_ ( .D(n7650), .CK(clock), .Q(
        decode_regfile_fpregs_13__16_) );
  DFF_X2 decode_regfile_fpregs_reg_13__17_ ( .D(n7649), .CK(clock), .Q(
        decode_regfile_fpregs_13__17_) );
  DFF_X2 decode_regfile_fpregs_reg_13__18_ ( .D(n7648), .CK(clock), .Q(
        decode_regfile_fpregs_13__18_) );
  DFF_X2 decode_regfile_fpregs_reg_13__19_ ( .D(n7647), .CK(clock), .Q(
        decode_regfile_fpregs_13__19_) );
  DFF_X2 decode_regfile_fpregs_reg_13__20_ ( .D(n7646), .CK(clock), .Q(
        decode_regfile_fpregs_13__20_) );
  DFF_X2 decode_regfile_fpregs_reg_13__21_ ( .D(n7645), .CK(clock), .Q(
        decode_regfile_fpregs_13__21_) );
  DFF_X2 decode_regfile_fpregs_reg_13__22_ ( .D(n7644), .CK(clock), .Q(
        decode_regfile_fpregs_13__22_) );
  DFF_X2 decode_regfile_fpregs_reg_13__23_ ( .D(n7643), .CK(clock), .Q(
        decode_regfile_fpregs_13__23_) );
  DFF_X2 decode_regfile_fpregs_reg_13__24_ ( .D(n7642), .CK(clock), .Q(
        decode_regfile_fpregs_13__24_) );
  DFF_X2 decode_regfile_fpregs_reg_13__25_ ( .D(n7641), .CK(clock), .Q(
        decode_regfile_fpregs_13__25_) );
  DFF_X2 decode_regfile_fpregs_reg_13__26_ ( .D(n7640), .CK(clock), .Q(
        decode_regfile_fpregs_13__26_) );
  DFF_X2 decode_regfile_fpregs_reg_13__27_ ( .D(n7639), .CK(clock), .Q(
        decode_regfile_fpregs_13__27_) );
  DFF_X2 decode_regfile_fpregs_reg_13__28_ ( .D(n7638), .CK(clock), .Q(
        decode_regfile_fpregs_13__28_) );
  DFF_X2 decode_regfile_fpregs_reg_13__29_ ( .D(n7637), .CK(clock), .Q(
        decode_regfile_fpregs_13__29_) );
  DFF_X2 decode_regfile_fpregs_reg_13__30_ ( .D(n7636), .CK(clock), .Q(
        decode_regfile_fpregs_13__30_) );
  DFF_X2 decode_regfile_fpregs_reg_13__31_ ( .D(n7635), .CK(clock), .Q(
        decode_regfile_fpregs_13__31_) );
  DFF_X2 decode_regfile_fpregs_reg_12__0_ ( .D(n7634), .CK(clock), .Q(
        decode_regfile_fpregs_12__0_) );
  DFF_X2 decode_regfile_fpregs_reg_12__1_ ( .D(n7633), .CK(clock), .Q(
        decode_regfile_fpregs_12__1_) );
  DFF_X2 decode_regfile_fpregs_reg_12__2_ ( .D(n7632), .CK(clock), .Q(
        decode_regfile_fpregs_12__2_) );
  DFF_X2 decode_regfile_fpregs_reg_12__3_ ( .D(n7631), .CK(clock), .Q(
        decode_regfile_fpregs_12__3_) );
  DFF_X2 decode_regfile_fpregs_reg_12__4_ ( .D(n7630), .CK(clock), .Q(
        decode_regfile_fpregs_12__4_) );
  DFF_X2 decode_regfile_fpregs_reg_12__5_ ( .D(n7629), .CK(clock), .Q(
        decode_regfile_fpregs_12__5_) );
  DFF_X2 decode_regfile_fpregs_reg_12__6_ ( .D(n7628), .CK(clock), .Q(
        decode_regfile_fpregs_12__6_) );
  DFF_X2 decode_regfile_fpregs_reg_12__7_ ( .D(n7627), .CK(clock), .Q(
        decode_regfile_fpregs_12__7_) );
  DFF_X2 decode_regfile_fpregs_reg_12__8_ ( .D(n7626), .CK(clock), .Q(
        decode_regfile_fpregs_12__8_) );
  DFF_X2 decode_regfile_fpregs_reg_12__9_ ( .D(n7625), .CK(clock), .Q(
        decode_regfile_fpregs_12__9_) );
  DFF_X2 decode_regfile_fpregs_reg_12__10_ ( .D(n7624), .CK(clock), .Q(
        decode_regfile_fpregs_12__10_) );
  DFF_X2 decode_regfile_fpregs_reg_12__11_ ( .D(n7623), .CK(clock), .Q(
        decode_regfile_fpregs_12__11_) );
  DFF_X2 decode_regfile_fpregs_reg_12__12_ ( .D(n7622), .CK(clock), .Q(
        decode_regfile_fpregs_12__12_) );
  DFF_X2 decode_regfile_fpregs_reg_12__13_ ( .D(n7621), .CK(clock), .Q(
        decode_regfile_fpregs_12__13_) );
  DFF_X2 decode_regfile_fpregs_reg_12__14_ ( .D(n7620), .CK(clock), .Q(
        decode_regfile_fpregs_12__14_) );
  DFF_X2 decode_regfile_fpregs_reg_12__15_ ( .D(n7619), .CK(clock), .Q(
        decode_regfile_fpregs_12__15_) );
  DFF_X2 decode_regfile_fpregs_reg_12__16_ ( .D(n7618), .CK(clock), .Q(
        decode_regfile_fpregs_12__16_) );
  DFF_X2 decode_regfile_fpregs_reg_12__17_ ( .D(n7617), .CK(clock), .Q(
        decode_regfile_fpregs_12__17_) );
  DFF_X2 decode_regfile_fpregs_reg_12__18_ ( .D(n7616), .CK(clock), .Q(
        decode_regfile_fpregs_12__18_) );
  DFF_X2 decode_regfile_fpregs_reg_12__19_ ( .D(n7615), .CK(clock), .Q(
        decode_regfile_fpregs_12__19_) );
  DFF_X2 decode_regfile_fpregs_reg_12__20_ ( .D(n7614), .CK(clock), .Q(
        decode_regfile_fpregs_12__20_) );
  DFF_X2 decode_regfile_fpregs_reg_12__21_ ( .D(n7613), .CK(clock), .Q(
        decode_regfile_fpregs_12__21_) );
  DFF_X2 decode_regfile_fpregs_reg_12__22_ ( .D(n7612), .CK(clock), .Q(
        decode_regfile_fpregs_12__22_) );
  DFF_X2 decode_regfile_fpregs_reg_12__23_ ( .D(n7611), .CK(clock), .Q(
        decode_regfile_fpregs_12__23_) );
  DFF_X2 decode_regfile_fpregs_reg_12__24_ ( .D(n7610), .CK(clock), .Q(
        decode_regfile_fpregs_12__24_) );
  DFF_X2 decode_regfile_fpregs_reg_12__25_ ( .D(n7609), .CK(clock), .Q(
        decode_regfile_fpregs_12__25_) );
  DFF_X2 decode_regfile_fpregs_reg_12__26_ ( .D(n7608), .CK(clock), .Q(
        decode_regfile_fpregs_12__26_) );
  DFF_X2 decode_regfile_fpregs_reg_12__27_ ( .D(n7607), .CK(clock), .Q(
        decode_regfile_fpregs_12__27_) );
  DFF_X2 decode_regfile_fpregs_reg_12__28_ ( .D(n7606), .CK(clock), .Q(
        decode_regfile_fpregs_12__28_) );
  DFF_X2 decode_regfile_fpregs_reg_12__29_ ( .D(n7605), .CK(clock), .Q(
        decode_regfile_fpregs_12__29_) );
  DFF_X2 decode_regfile_fpregs_reg_12__30_ ( .D(n7604), .CK(clock), .Q(
        decode_regfile_fpregs_12__30_) );
  DFF_X2 decode_regfile_fpregs_reg_12__31_ ( .D(n7603), .CK(clock), .Q(
        decode_regfile_fpregs_12__31_) );
  DFF_X2 decode_regfile_fpregs_reg_11__0_ ( .D(n7602), .CK(clock), .Q(
        decode_regfile_fpregs_11__0_) );
  DFF_X2 decode_regfile_fpregs_reg_11__1_ ( .D(n7601), .CK(clock), .Q(
        decode_regfile_fpregs_11__1_) );
  DFF_X2 decode_regfile_fpregs_reg_11__2_ ( .D(n7600), .CK(clock), .Q(
        decode_regfile_fpregs_11__2_) );
  DFF_X2 decode_regfile_fpregs_reg_11__3_ ( .D(n7599), .CK(clock), .Q(
        decode_regfile_fpregs_11__3_) );
  DFF_X2 decode_regfile_fpregs_reg_11__4_ ( .D(n7598), .CK(clock), .Q(
        decode_regfile_fpregs_11__4_) );
  DFF_X2 decode_regfile_fpregs_reg_11__5_ ( .D(n7597), .CK(clock), .Q(
        decode_regfile_fpregs_11__5_) );
  DFF_X2 decode_regfile_fpregs_reg_11__6_ ( .D(n7596), .CK(clock), .Q(
        decode_regfile_fpregs_11__6_) );
  DFF_X2 decode_regfile_fpregs_reg_11__7_ ( .D(n7595), .CK(clock), .Q(
        decode_regfile_fpregs_11__7_) );
  DFF_X2 decode_regfile_fpregs_reg_11__8_ ( .D(n7594), .CK(clock), .Q(
        decode_regfile_fpregs_11__8_) );
  DFF_X2 decode_regfile_fpregs_reg_11__9_ ( .D(n7593), .CK(clock), .Q(
        decode_regfile_fpregs_11__9_) );
  DFF_X2 decode_regfile_fpregs_reg_11__10_ ( .D(n7592), .CK(clock), .Q(
        decode_regfile_fpregs_11__10_) );
  DFF_X2 decode_regfile_fpregs_reg_11__11_ ( .D(n7591), .CK(clock), .Q(
        decode_regfile_fpregs_11__11_) );
  DFF_X2 decode_regfile_fpregs_reg_11__12_ ( .D(n7590), .CK(clock), .Q(
        decode_regfile_fpregs_11__12_) );
  DFF_X2 decode_regfile_fpregs_reg_11__13_ ( .D(n7589), .CK(clock), .Q(
        decode_regfile_fpregs_11__13_) );
  DFF_X2 decode_regfile_fpregs_reg_11__14_ ( .D(n7588), .CK(clock), .Q(
        decode_regfile_fpregs_11__14_) );
  DFF_X2 decode_regfile_fpregs_reg_11__15_ ( .D(n7587), .CK(clock), .Q(
        decode_regfile_fpregs_11__15_) );
  DFF_X2 decode_regfile_fpregs_reg_11__16_ ( .D(n7586), .CK(clock), .Q(
        decode_regfile_fpregs_11__16_) );
  DFF_X2 decode_regfile_fpregs_reg_11__17_ ( .D(n7585), .CK(clock), .Q(
        decode_regfile_fpregs_11__17_) );
  DFF_X2 decode_regfile_fpregs_reg_11__18_ ( .D(n7584), .CK(clock), .Q(
        decode_regfile_fpregs_11__18_) );
  DFF_X2 decode_regfile_fpregs_reg_11__19_ ( .D(n7583), .CK(clock), .Q(
        decode_regfile_fpregs_11__19_) );
  DFF_X2 decode_regfile_fpregs_reg_11__20_ ( .D(n7582), .CK(clock), .Q(
        decode_regfile_fpregs_11__20_) );
  DFF_X2 decode_regfile_fpregs_reg_11__21_ ( .D(n7581), .CK(clock), .Q(
        decode_regfile_fpregs_11__21_) );
  DFF_X2 decode_regfile_fpregs_reg_11__22_ ( .D(n7580), .CK(clock), .Q(
        decode_regfile_fpregs_11__22_) );
  DFF_X2 decode_regfile_fpregs_reg_11__23_ ( .D(n7579), .CK(clock), .Q(
        decode_regfile_fpregs_11__23_) );
  DFF_X2 decode_regfile_fpregs_reg_11__24_ ( .D(n7578), .CK(clock), .Q(
        decode_regfile_fpregs_11__24_) );
  DFF_X2 decode_regfile_fpregs_reg_11__25_ ( .D(n7577), .CK(clock), .Q(
        decode_regfile_fpregs_11__25_) );
  DFF_X2 decode_regfile_fpregs_reg_11__26_ ( .D(n7576), .CK(clock), .Q(
        decode_regfile_fpregs_11__26_) );
  DFF_X2 decode_regfile_fpregs_reg_11__27_ ( .D(n7575), .CK(clock), .Q(
        decode_regfile_fpregs_11__27_) );
  DFF_X2 decode_regfile_fpregs_reg_11__28_ ( .D(n7574), .CK(clock), .Q(
        decode_regfile_fpregs_11__28_) );
  DFF_X2 decode_regfile_fpregs_reg_11__29_ ( .D(n7573), .CK(clock), .Q(
        decode_regfile_fpregs_11__29_) );
  DFF_X2 decode_regfile_fpregs_reg_11__30_ ( .D(n7572), .CK(clock), .Q(
        decode_regfile_fpregs_11__30_) );
  DFF_X2 decode_regfile_fpregs_reg_11__31_ ( .D(n7571), .CK(clock), .Q(
        decode_regfile_fpregs_11__31_) );
  DFF_X2 decode_regfile_fpregs_reg_10__0_ ( .D(n7570), .CK(clock), .Q(
        decode_regfile_fpregs_10__0_) );
  DFF_X2 decode_regfile_fpregs_reg_10__1_ ( .D(n7569), .CK(clock), .Q(
        decode_regfile_fpregs_10__1_) );
  DFF_X2 decode_regfile_fpregs_reg_10__2_ ( .D(n7568), .CK(clock), .Q(
        decode_regfile_fpregs_10__2_) );
  DFF_X2 decode_regfile_fpregs_reg_10__3_ ( .D(n7567), .CK(clock), .Q(
        decode_regfile_fpregs_10__3_) );
  DFF_X2 decode_regfile_fpregs_reg_10__4_ ( .D(n7566), .CK(clock), .Q(
        decode_regfile_fpregs_10__4_) );
  DFF_X2 decode_regfile_fpregs_reg_10__5_ ( .D(n7565), .CK(clock), .Q(
        decode_regfile_fpregs_10__5_) );
  DFF_X2 decode_regfile_fpregs_reg_10__6_ ( .D(n7564), .CK(clock), .Q(
        decode_regfile_fpregs_10__6_) );
  DFF_X2 decode_regfile_fpregs_reg_10__7_ ( .D(n7563), .CK(clock), .Q(
        decode_regfile_fpregs_10__7_) );
  DFF_X2 decode_regfile_fpregs_reg_10__8_ ( .D(n7562), .CK(clock), .Q(
        decode_regfile_fpregs_10__8_) );
  DFF_X2 decode_regfile_fpregs_reg_10__9_ ( .D(n7561), .CK(clock), .Q(
        decode_regfile_fpregs_10__9_) );
  DFF_X2 decode_regfile_fpregs_reg_10__10_ ( .D(n7560), .CK(clock), .Q(
        decode_regfile_fpregs_10__10_) );
  DFF_X2 decode_regfile_fpregs_reg_10__11_ ( .D(n7559), .CK(clock), .Q(
        decode_regfile_fpregs_10__11_) );
  DFF_X2 decode_regfile_fpregs_reg_10__12_ ( .D(n7558), .CK(clock), .Q(
        decode_regfile_fpregs_10__12_) );
  DFF_X2 decode_regfile_fpregs_reg_10__13_ ( .D(n7557), .CK(clock), .Q(
        decode_regfile_fpregs_10__13_) );
  DFF_X2 decode_regfile_fpregs_reg_10__14_ ( .D(n7556), .CK(clock), .Q(
        decode_regfile_fpregs_10__14_) );
  DFF_X2 decode_regfile_fpregs_reg_10__15_ ( .D(n7555), .CK(clock), .Q(
        decode_regfile_fpregs_10__15_) );
  DFF_X2 decode_regfile_fpregs_reg_10__16_ ( .D(n7554), .CK(clock), .Q(
        decode_regfile_fpregs_10__16_) );
  DFF_X2 decode_regfile_fpregs_reg_10__17_ ( .D(n7553), .CK(clock), .Q(
        decode_regfile_fpregs_10__17_) );
  DFF_X2 decode_regfile_fpregs_reg_10__18_ ( .D(n7552), .CK(clock), .Q(
        decode_regfile_fpregs_10__18_) );
  DFF_X2 decode_regfile_fpregs_reg_10__19_ ( .D(n7551), .CK(clock), .Q(
        decode_regfile_fpregs_10__19_) );
  DFF_X2 decode_regfile_fpregs_reg_10__20_ ( .D(n7550), .CK(clock), .Q(
        decode_regfile_fpregs_10__20_) );
  DFF_X2 decode_regfile_fpregs_reg_10__21_ ( .D(n7549), .CK(clock), .Q(
        decode_regfile_fpregs_10__21_) );
  DFF_X2 decode_regfile_fpregs_reg_10__22_ ( .D(n7548), .CK(clock), .Q(
        decode_regfile_fpregs_10__22_) );
  DFF_X2 decode_regfile_fpregs_reg_10__23_ ( .D(n7547), .CK(clock), .Q(
        decode_regfile_fpregs_10__23_) );
  DFF_X2 decode_regfile_fpregs_reg_10__24_ ( .D(n7546), .CK(clock), .Q(
        decode_regfile_fpregs_10__24_) );
  DFF_X2 decode_regfile_fpregs_reg_10__25_ ( .D(n7545), .CK(clock), .Q(
        decode_regfile_fpregs_10__25_) );
  DFF_X2 decode_regfile_fpregs_reg_10__26_ ( .D(n7544), .CK(clock), .Q(
        decode_regfile_fpregs_10__26_) );
  DFF_X2 decode_regfile_fpregs_reg_10__27_ ( .D(n7543), .CK(clock), .Q(
        decode_regfile_fpregs_10__27_) );
  DFF_X2 decode_regfile_fpregs_reg_10__28_ ( .D(n7542), .CK(clock), .Q(
        decode_regfile_fpregs_10__28_) );
  DFF_X2 decode_regfile_fpregs_reg_10__29_ ( .D(n7541), .CK(clock), .Q(
        decode_regfile_fpregs_10__29_) );
  DFF_X2 decode_regfile_fpregs_reg_10__30_ ( .D(n7540), .CK(clock), .Q(
        decode_regfile_fpregs_10__30_) );
  DFF_X2 decode_regfile_fpregs_reg_10__31_ ( .D(n7539), .CK(clock), .Q(
        decode_regfile_fpregs_10__31_) );
  DFF_X2 decode_regfile_fpregs_reg_9__0_ ( .D(n7538), .CK(clock), .Q(
        decode_regfile_fpregs_9__0_) );
  DFF_X2 decode_regfile_fpregs_reg_9__1_ ( .D(n7537), .CK(clock), .Q(
        decode_regfile_fpregs_9__1_) );
  DFF_X2 decode_regfile_fpregs_reg_9__2_ ( .D(n7536), .CK(clock), .Q(
        decode_regfile_fpregs_9__2_) );
  DFF_X2 decode_regfile_fpregs_reg_9__3_ ( .D(n7535), .CK(clock), .Q(
        decode_regfile_fpregs_9__3_) );
  DFF_X2 decode_regfile_fpregs_reg_9__4_ ( .D(n7534), .CK(clock), .Q(
        decode_regfile_fpregs_9__4_) );
  DFF_X2 decode_regfile_fpregs_reg_9__5_ ( .D(n7533), .CK(clock), .Q(
        decode_regfile_fpregs_9__5_) );
  DFF_X2 decode_regfile_fpregs_reg_9__6_ ( .D(n7532), .CK(clock), .Q(
        decode_regfile_fpregs_9__6_) );
  DFF_X2 decode_regfile_fpregs_reg_9__7_ ( .D(n7531), .CK(clock), .Q(
        decode_regfile_fpregs_9__7_) );
  DFF_X2 decode_regfile_fpregs_reg_9__8_ ( .D(n7530), .CK(clock), .Q(
        decode_regfile_fpregs_9__8_) );
  DFF_X2 decode_regfile_fpregs_reg_9__9_ ( .D(n7529), .CK(clock), .Q(
        decode_regfile_fpregs_9__9_) );
  DFF_X2 decode_regfile_fpregs_reg_9__10_ ( .D(n7528), .CK(clock), .Q(
        decode_regfile_fpregs_9__10_) );
  DFF_X2 decode_regfile_fpregs_reg_9__11_ ( .D(n7527), .CK(clock), .Q(
        decode_regfile_fpregs_9__11_) );
  DFF_X2 decode_regfile_fpregs_reg_9__12_ ( .D(n7526), .CK(clock), .Q(
        decode_regfile_fpregs_9__12_) );
  DFF_X2 decode_regfile_fpregs_reg_9__13_ ( .D(n7525), .CK(clock), .Q(
        decode_regfile_fpregs_9__13_) );
  DFF_X2 decode_regfile_fpregs_reg_9__14_ ( .D(n7524), .CK(clock), .Q(
        decode_regfile_fpregs_9__14_) );
  DFF_X2 decode_regfile_fpregs_reg_9__15_ ( .D(n7523), .CK(clock), .Q(
        decode_regfile_fpregs_9__15_) );
  DFF_X2 decode_regfile_fpregs_reg_9__16_ ( .D(n7522), .CK(clock), .Q(
        decode_regfile_fpregs_9__16_) );
  DFF_X2 decode_regfile_fpregs_reg_9__17_ ( .D(n7521), .CK(clock), .Q(
        decode_regfile_fpregs_9__17_) );
  DFF_X2 decode_regfile_fpregs_reg_9__18_ ( .D(n7520), .CK(clock), .Q(
        decode_regfile_fpregs_9__18_) );
  DFF_X2 decode_regfile_fpregs_reg_9__19_ ( .D(n7519), .CK(clock), .Q(
        decode_regfile_fpregs_9__19_) );
  DFF_X2 decode_regfile_fpregs_reg_9__20_ ( .D(n7518), .CK(clock), .Q(
        decode_regfile_fpregs_9__20_) );
  DFF_X2 decode_regfile_fpregs_reg_9__21_ ( .D(n7517), .CK(clock), .Q(
        decode_regfile_fpregs_9__21_) );
  DFF_X2 decode_regfile_fpregs_reg_9__22_ ( .D(n7516), .CK(clock), .Q(
        decode_regfile_fpregs_9__22_) );
  DFF_X2 decode_regfile_fpregs_reg_9__23_ ( .D(n7515), .CK(clock), .Q(
        decode_regfile_fpregs_9__23_) );
  DFF_X2 decode_regfile_fpregs_reg_9__24_ ( .D(n7514), .CK(clock), .Q(
        decode_regfile_fpregs_9__24_) );
  DFF_X2 decode_regfile_fpregs_reg_9__25_ ( .D(n7513), .CK(clock), .Q(
        decode_regfile_fpregs_9__25_) );
  DFF_X2 decode_regfile_fpregs_reg_9__26_ ( .D(n7512), .CK(clock), .Q(
        decode_regfile_fpregs_9__26_) );
  DFF_X2 decode_regfile_fpregs_reg_9__27_ ( .D(n7511), .CK(clock), .Q(
        decode_regfile_fpregs_9__27_) );
  DFF_X2 decode_regfile_fpregs_reg_9__28_ ( .D(n7510), .CK(clock), .Q(
        decode_regfile_fpregs_9__28_) );
  DFF_X2 decode_regfile_fpregs_reg_9__29_ ( .D(n7509), .CK(clock), .Q(
        decode_regfile_fpregs_9__29_) );
  DFF_X2 decode_regfile_fpregs_reg_9__30_ ( .D(n7508), .CK(clock), .Q(
        decode_regfile_fpregs_9__30_) );
  DFF_X2 decode_regfile_fpregs_reg_9__31_ ( .D(n7507), .CK(clock), .Q(
        decode_regfile_fpregs_9__31_) );
  DFF_X2 decode_regfile_fpregs_reg_8__0_ ( .D(n7506), .CK(clock), .Q(
        decode_regfile_fpregs_8__0_) );
  DFF_X2 decode_regfile_fpregs_reg_8__1_ ( .D(n7505), .CK(clock), .Q(
        decode_regfile_fpregs_8__1_) );
  DFF_X2 decode_regfile_fpregs_reg_8__2_ ( .D(n7504), .CK(clock), .Q(
        decode_regfile_fpregs_8__2_) );
  DFF_X2 decode_regfile_fpregs_reg_8__3_ ( .D(n7503), .CK(clock), .Q(
        decode_regfile_fpregs_8__3_) );
  DFF_X2 decode_regfile_fpregs_reg_8__4_ ( .D(n7502), .CK(clock), .Q(
        decode_regfile_fpregs_8__4_) );
  DFF_X2 decode_regfile_fpregs_reg_8__5_ ( .D(n7501), .CK(clock), .Q(
        decode_regfile_fpregs_8__5_) );
  DFF_X2 decode_regfile_fpregs_reg_8__6_ ( .D(n7500), .CK(clock), .Q(
        decode_regfile_fpregs_8__6_) );
  DFF_X2 decode_regfile_fpregs_reg_8__7_ ( .D(n7499), .CK(clock), .Q(
        decode_regfile_fpregs_8__7_) );
  DFF_X2 decode_regfile_fpregs_reg_8__8_ ( .D(n7498), .CK(clock), .Q(
        decode_regfile_fpregs_8__8_) );
  DFF_X2 decode_regfile_fpregs_reg_8__9_ ( .D(n7497), .CK(clock), .Q(
        decode_regfile_fpregs_8__9_) );
  DFF_X2 decode_regfile_fpregs_reg_8__10_ ( .D(n7496), .CK(clock), .Q(
        decode_regfile_fpregs_8__10_) );
  DFF_X2 decode_regfile_fpregs_reg_8__11_ ( .D(n7495), .CK(clock), .Q(
        decode_regfile_fpregs_8__11_) );
  DFF_X2 decode_regfile_fpregs_reg_8__12_ ( .D(n7494), .CK(clock), .Q(
        decode_regfile_fpregs_8__12_) );
  DFF_X2 decode_regfile_fpregs_reg_8__13_ ( .D(n7493), .CK(clock), .Q(
        decode_regfile_fpregs_8__13_) );
  DFF_X2 decode_regfile_fpregs_reg_8__14_ ( .D(n7492), .CK(clock), .Q(
        decode_regfile_fpregs_8__14_) );
  DFF_X2 decode_regfile_fpregs_reg_8__15_ ( .D(n7491), .CK(clock), .Q(
        decode_regfile_fpregs_8__15_) );
  DFF_X2 decode_regfile_fpregs_reg_8__16_ ( .D(n7490), .CK(clock), .Q(
        decode_regfile_fpregs_8__16_) );
  DFF_X2 decode_regfile_fpregs_reg_8__17_ ( .D(n7489), .CK(clock), .Q(
        decode_regfile_fpregs_8__17_) );
  DFF_X2 decode_regfile_fpregs_reg_8__18_ ( .D(n7488), .CK(clock), .Q(
        decode_regfile_fpregs_8__18_) );
  DFF_X2 decode_regfile_fpregs_reg_8__19_ ( .D(n7487), .CK(clock), .Q(
        decode_regfile_fpregs_8__19_) );
  DFF_X2 decode_regfile_fpregs_reg_8__20_ ( .D(n7486), .CK(clock), .Q(
        decode_regfile_fpregs_8__20_) );
  DFF_X2 decode_regfile_fpregs_reg_8__21_ ( .D(n7485), .CK(clock), .Q(
        decode_regfile_fpregs_8__21_) );
  DFF_X2 decode_regfile_fpregs_reg_8__22_ ( .D(n7484), .CK(clock), .Q(
        decode_regfile_fpregs_8__22_) );
  DFF_X2 decode_regfile_fpregs_reg_8__23_ ( .D(n7483), .CK(clock), .Q(
        decode_regfile_fpregs_8__23_) );
  DFF_X2 decode_regfile_fpregs_reg_8__24_ ( .D(n7482), .CK(clock), .Q(
        decode_regfile_fpregs_8__24_) );
  DFF_X2 decode_regfile_fpregs_reg_8__25_ ( .D(n7481), .CK(clock), .Q(
        decode_regfile_fpregs_8__25_) );
  DFF_X2 decode_regfile_fpregs_reg_8__26_ ( .D(n7480), .CK(clock), .Q(
        decode_regfile_fpregs_8__26_) );
  DFF_X2 decode_regfile_fpregs_reg_8__27_ ( .D(n7479), .CK(clock), .Q(
        decode_regfile_fpregs_8__27_) );
  DFF_X2 decode_regfile_fpregs_reg_8__28_ ( .D(n7478), .CK(clock), .Q(
        decode_regfile_fpregs_8__28_) );
  DFF_X2 decode_regfile_fpregs_reg_8__29_ ( .D(n7477), .CK(clock), .Q(
        decode_regfile_fpregs_8__29_) );
  DFF_X2 decode_regfile_fpregs_reg_8__30_ ( .D(n7476), .CK(clock), .Q(
        decode_regfile_fpregs_8__30_) );
  DFF_X2 decode_regfile_fpregs_reg_8__31_ ( .D(n7475), .CK(clock), .Q(
        decode_regfile_fpregs_8__31_) );
  DFF_X2 decode_regfile_fpregs_reg_7__0_ ( .D(n7474), .CK(clock), .Q(
        decode_regfile_fpregs_7__0_) );
  DFF_X2 decode_regfile_fpregs_reg_7__1_ ( .D(n7473), .CK(clock), .Q(
        decode_regfile_fpregs_7__1_) );
  DFF_X2 decode_regfile_fpregs_reg_7__2_ ( .D(n7472), .CK(clock), .Q(
        decode_regfile_fpregs_7__2_) );
  DFF_X2 decode_regfile_fpregs_reg_7__3_ ( .D(n7471), .CK(clock), .Q(
        decode_regfile_fpregs_7__3_) );
  DFF_X2 decode_regfile_fpregs_reg_7__4_ ( .D(n7470), .CK(clock), .Q(
        decode_regfile_fpregs_7__4_) );
  DFF_X2 decode_regfile_fpregs_reg_7__5_ ( .D(n7469), .CK(clock), .Q(
        decode_regfile_fpregs_7__5_) );
  DFF_X2 decode_regfile_fpregs_reg_7__6_ ( .D(n7468), .CK(clock), .Q(
        decode_regfile_fpregs_7__6_) );
  DFF_X2 decode_regfile_fpregs_reg_7__7_ ( .D(n7467), .CK(clock), .Q(
        decode_regfile_fpregs_7__7_) );
  DFF_X2 decode_regfile_fpregs_reg_7__8_ ( .D(n7466), .CK(clock), .Q(
        decode_regfile_fpregs_7__8_) );
  DFF_X2 decode_regfile_fpregs_reg_7__9_ ( .D(n7465), .CK(clock), .Q(
        decode_regfile_fpregs_7__9_) );
  DFF_X2 decode_regfile_fpregs_reg_7__10_ ( .D(n7464), .CK(clock), .Q(
        decode_regfile_fpregs_7__10_) );
  DFF_X2 decode_regfile_fpregs_reg_7__11_ ( .D(n7463), .CK(clock), .Q(
        decode_regfile_fpregs_7__11_) );
  DFF_X2 decode_regfile_fpregs_reg_7__12_ ( .D(n7462), .CK(clock), .Q(
        decode_regfile_fpregs_7__12_) );
  DFF_X2 decode_regfile_fpregs_reg_7__13_ ( .D(n7461), .CK(clock), .Q(
        decode_regfile_fpregs_7__13_) );
  DFF_X2 decode_regfile_fpregs_reg_7__14_ ( .D(n7460), .CK(clock), .Q(
        decode_regfile_fpregs_7__14_) );
  DFF_X2 decode_regfile_fpregs_reg_7__15_ ( .D(n7459), .CK(clock), .Q(
        decode_regfile_fpregs_7__15_) );
  DFF_X2 decode_regfile_fpregs_reg_7__16_ ( .D(n7458), .CK(clock), .Q(
        decode_regfile_fpregs_7__16_) );
  DFF_X2 decode_regfile_fpregs_reg_7__17_ ( .D(n7457), .CK(clock), .Q(
        decode_regfile_fpregs_7__17_) );
  DFF_X2 decode_regfile_fpregs_reg_7__18_ ( .D(n7456), .CK(clock), .Q(
        decode_regfile_fpregs_7__18_) );
  DFF_X2 decode_regfile_fpregs_reg_7__19_ ( .D(n7455), .CK(clock), .Q(
        decode_regfile_fpregs_7__19_) );
  DFF_X2 decode_regfile_fpregs_reg_7__20_ ( .D(n7454), .CK(clock), .Q(
        decode_regfile_fpregs_7__20_) );
  DFF_X2 decode_regfile_fpregs_reg_7__21_ ( .D(n7453), .CK(clock), .Q(
        decode_regfile_fpregs_7__21_) );
  DFF_X2 decode_regfile_fpregs_reg_7__22_ ( .D(n7452), .CK(clock), .Q(
        decode_regfile_fpregs_7__22_) );
  DFF_X2 decode_regfile_fpregs_reg_7__23_ ( .D(n7451), .CK(clock), .Q(
        decode_regfile_fpregs_7__23_) );
  DFF_X2 decode_regfile_fpregs_reg_7__24_ ( .D(n7450), .CK(clock), .Q(
        decode_regfile_fpregs_7__24_) );
  DFF_X2 decode_regfile_fpregs_reg_7__25_ ( .D(n7449), .CK(clock), .Q(
        decode_regfile_fpregs_7__25_) );
  DFF_X2 decode_regfile_fpregs_reg_7__26_ ( .D(n7448), .CK(clock), .Q(
        decode_regfile_fpregs_7__26_) );
  DFF_X2 decode_regfile_fpregs_reg_7__27_ ( .D(n7447), .CK(clock), .Q(
        decode_regfile_fpregs_7__27_) );
  DFF_X2 decode_regfile_fpregs_reg_7__28_ ( .D(n7446), .CK(clock), .Q(
        decode_regfile_fpregs_7__28_) );
  DFF_X2 decode_regfile_fpregs_reg_7__29_ ( .D(n7445), .CK(clock), .Q(
        decode_regfile_fpregs_7__29_) );
  DFF_X2 decode_regfile_fpregs_reg_7__30_ ( .D(n7444), .CK(clock), .Q(
        decode_regfile_fpregs_7__30_) );
  DFF_X2 decode_regfile_fpregs_reg_7__31_ ( .D(n7443), .CK(clock), .Q(
        decode_regfile_fpregs_7__31_) );
  DFF_X2 decode_regfile_fpregs_reg_6__0_ ( .D(n7442), .CK(clock), .Q(
        decode_regfile_fpregs_6__0_) );
  DFF_X2 decode_regfile_fpregs_reg_6__1_ ( .D(n7441), .CK(clock), .Q(
        decode_regfile_fpregs_6__1_) );
  DFF_X2 decode_regfile_fpregs_reg_6__2_ ( .D(n7440), .CK(clock), .Q(
        decode_regfile_fpregs_6__2_) );
  DFF_X2 decode_regfile_fpregs_reg_6__3_ ( .D(n7439), .CK(clock), .Q(
        decode_regfile_fpregs_6__3_) );
  DFF_X2 decode_regfile_fpregs_reg_6__4_ ( .D(n7438), .CK(clock), .Q(
        decode_regfile_fpregs_6__4_) );
  DFF_X2 decode_regfile_fpregs_reg_6__5_ ( .D(n7437), .CK(clock), .Q(
        decode_regfile_fpregs_6__5_) );
  DFF_X2 decode_regfile_fpregs_reg_6__6_ ( .D(n7436), .CK(clock), .Q(
        decode_regfile_fpregs_6__6_) );
  DFF_X2 decode_regfile_fpregs_reg_6__7_ ( .D(n7435), .CK(clock), .Q(
        decode_regfile_fpregs_6__7_) );
  DFF_X2 decode_regfile_fpregs_reg_6__8_ ( .D(n7434), .CK(clock), .Q(
        decode_regfile_fpregs_6__8_) );
  DFF_X2 decode_regfile_fpregs_reg_6__9_ ( .D(n7433), .CK(clock), .Q(
        decode_regfile_fpregs_6__9_) );
  DFF_X2 decode_regfile_fpregs_reg_6__10_ ( .D(n7432), .CK(clock), .Q(
        decode_regfile_fpregs_6__10_) );
  DFF_X2 decode_regfile_fpregs_reg_6__11_ ( .D(n7431), .CK(clock), .Q(
        decode_regfile_fpregs_6__11_) );
  DFF_X2 decode_regfile_fpregs_reg_6__12_ ( .D(n7430), .CK(clock), .Q(
        decode_regfile_fpregs_6__12_) );
  DFF_X2 decode_regfile_fpregs_reg_6__13_ ( .D(n7429), .CK(clock), .Q(
        decode_regfile_fpregs_6__13_) );
  DFF_X2 decode_regfile_fpregs_reg_6__14_ ( .D(n7428), .CK(clock), .Q(
        decode_regfile_fpregs_6__14_) );
  DFF_X2 decode_regfile_fpregs_reg_6__15_ ( .D(n7427), .CK(clock), .Q(
        decode_regfile_fpregs_6__15_) );
  DFF_X2 decode_regfile_fpregs_reg_6__16_ ( .D(n7426), .CK(clock), .Q(
        decode_regfile_fpregs_6__16_) );
  DFF_X2 decode_regfile_fpregs_reg_6__17_ ( .D(n7425), .CK(clock), .Q(
        decode_regfile_fpregs_6__17_) );
  DFF_X2 decode_regfile_fpregs_reg_6__18_ ( .D(n7424), .CK(clock), .Q(
        decode_regfile_fpregs_6__18_) );
  DFF_X2 decode_regfile_fpregs_reg_6__19_ ( .D(n7423), .CK(clock), .Q(
        decode_regfile_fpregs_6__19_) );
  DFF_X2 decode_regfile_fpregs_reg_6__20_ ( .D(n7422), .CK(clock), .Q(
        decode_regfile_fpregs_6__20_) );
  DFF_X2 decode_regfile_fpregs_reg_6__21_ ( .D(n7421), .CK(clock), .Q(
        decode_regfile_fpregs_6__21_) );
  DFF_X2 decode_regfile_fpregs_reg_6__22_ ( .D(n7420), .CK(clock), .Q(
        decode_regfile_fpregs_6__22_) );
  DFF_X2 decode_regfile_fpregs_reg_6__23_ ( .D(n7419), .CK(clock), .Q(
        decode_regfile_fpregs_6__23_) );
  DFF_X2 decode_regfile_fpregs_reg_6__24_ ( .D(n7418), .CK(clock), .Q(
        decode_regfile_fpregs_6__24_) );
  DFF_X2 decode_regfile_fpregs_reg_6__25_ ( .D(n7417), .CK(clock), .Q(
        decode_regfile_fpregs_6__25_) );
  DFF_X2 decode_regfile_fpregs_reg_6__26_ ( .D(n7416), .CK(clock), .Q(
        decode_regfile_fpregs_6__26_) );
  DFF_X2 decode_regfile_fpregs_reg_6__27_ ( .D(n7415), .CK(clock), .Q(
        decode_regfile_fpregs_6__27_) );
  DFF_X2 decode_regfile_fpregs_reg_6__28_ ( .D(n7414), .CK(clock), .Q(
        decode_regfile_fpregs_6__28_) );
  DFF_X2 decode_regfile_fpregs_reg_6__29_ ( .D(n7413), .CK(clock), .Q(
        decode_regfile_fpregs_6__29_) );
  DFF_X2 decode_regfile_fpregs_reg_6__30_ ( .D(n7412), .CK(clock), .Q(
        decode_regfile_fpregs_6__30_) );
  DFF_X2 decode_regfile_fpregs_reg_6__31_ ( .D(n7411), .CK(clock), .Q(
        decode_regfile_fpregs_6__31_) );
  DFF_X2 decode_regfile_fpregs_reg_5__0_ ( .D(n7410), .CK(clock), .Q(
        decode_regfile_fpregs_5__0_) );
  DFF_X2 decode_regfile_fpregs_reg_5__1_ ( .D(n7409), .CK(clock), .Q(
        decode_regfile_fpregs_5__1_) );
  DFF_X2 decode_regfile_fpregs_reg_5__2_ ( .D(n7408), .CK(clock), .Q(
        decode_regfile_fpregs_5__2_) );
  DFF_X2 decode_regfile_fpregs_reg_5__3_ ( .D(n7407), .CK(clock), .Q(
        decode_regfile_fpregs_5__3_) );
  DFF_X2 decode_regfile_fpregs_reg_5__4_ ( .D(n7406), .CK(clock), .Q(
        decode_regfile_fpregs_5__4_) );
  DFF_X2 decode_regfile_fpregs_reg_5__5_ ( .D(n7405), .CK(clock), .Q(
        decode_regfile_fpregs_5__5_) );
  DFF_X2 decode_regfile_fpregs_reg_5__6_ ( .D(n7404), .CK(clock), .Q(
        decode_regfile_fpregs_5__6_) );
  DFF_X2 decode_regfile_fpregs_reg_5__7_ ( .D(n7403), .CK(clock), .Q(
        decode_regfile_fpregs_5__7_) );
  DFF_X2 decode_regfile_fpregs_reg_5__8_ ( .D(n7402), .CK(clock), .Q(
        decode_regfile_fpregs_5__8_) );
  DFF_X2 decode_regfile_fpregs_reg_5__9_ ( .D(n7401), .CK(clock), .Q(
        decode_regfile_fpregs_5__9_) );
  DFF_X2 decode_regfile_fpregs_reg_5__10_ ( .D(n7400), .CK(clock), .Q(
        decode_regfile_fpregs_5__10_) );
  DFF_X2 decode_regfile_fpregs_reg_5__11_ ( .D(n7399), .CK(clock), .Q(
        decode_regfile_fpregs_5__11_) );
  DFF_X2 decode_regfile_fpregs_reg_5__12_ ( .D(n7398), .CK(clock), .Q(
        decode_regfile_fpregs_5__12_) );
  DFF_X2 decode_regfile_fpregs_reg_5__13_ ( .D(n7397), .CK(clock), .Q(
        decode_regfile_fpregs_5__13_) );
  DFF_X2 decode_regfile_fpregs_reg_5__14_ ( .D(n7396), .CK(clock), .Q(
        decode_regfile_fpregs_5__14_) );
  DFF_X2 decode_regfile_fpregs_reg_5__15_ ( .D(n7395), .CK(clock), .Q(
        decode_regfile_fpregs_5__15_) );
  DFF_X2 decode_regfile_fpregs_reg_5__16_ ( .D(n7394), .CK(clock), .Q(
        decode_regfile_fpregs_5__16_) );
  DFF_X2 decode_regfile_fpregs_reg_5__17_ ( .D(n7393), .CK(clock), .Q(
        decode_regfile_fpregs_5__17_) );
  DFF_X2 decode_regfile_fpregs_reg_5__18_ ( .D(n7392), .CK(clock), .Q(
        decode_regfile_fpregs_5__18_) );
  DFF_X2 decode_regfile_fpregs_reg_5__19_ ( .D(n7391), .CK(clock), .Q(
        decode_regfile_fpregs_5__19_) );
  DFF_X2 decode_regfile_fpregs_reg_5__20_ ( .D(n7390), .CK(clock), .Q(
        decode_regfile_fpregs_5__20_) );
  DFF_X2 decode_regfile_fpregs_reg_5__21_ ( .D(n7389), .CK(clock), .Q(
        decode_regfile_fpregs_5__21_) );
  DFF_X2 decode_regfile_fpregs_reg_5__22_ ( .D(n7388), .CK(clock), .Q(
        decode_regfile_fpregs_5__22_) );
  DFF_X2 decode_regfile_fpregs_reg_5__23_ ( .D(n7387), .CK(clock), .Q(
        decode_regfile_fpregs_5__23_) );
  DFF_X2 decode_regfile_fpregs_reg_5__24_ ( .D(n7386), .CK(clock), .Q(
        decode_regfile_fpregs_5__24_) );
  DFF_X2 decode_regfile_fpregs_reg_5__25_ ( .D(n7385), .CK(clock), .Q(
        decode_regfile_fpregs_5__25_) );
  DFF_X2 decode_regfile_fpregs_reg_5__26_ ( .D(n7384), .CK(clock), .Q(
        decode_regfile_fpregs_5__26_) );
  DFF_X2 decode_regfile_fpregs_reg_5__27_ ( .D(n7383), .CK(clock), .Q(
        decode_regfile_fpregs_5__27_) );
  DFF_X2 decode_regfile_fpregs_reg_5__28_ ( .D(n7382), .CK(clock), .Q(
        decode_regfile_fpregs_5__28_) );
  DFF_X2 decode_regfile_fpregs_reg_5__29_ ( .D(n7381), .CK(clock), .Q(
        decode_regfile_fpregs_5__29_) );
  DFF_X2 decode_regfile_fpregs_reg_5__30_ ( .D(n7380), .CK(clock), .Q(
        decode_regfile_fpregs_5__30_) );
  DFF_X2 decode_regfile_fpregs_reg_5__31_ ( .D(n7379), .CK(clock), .Q(
        decode_regfile_fpregs_5__31_) );
  DFF_X2 decode_regfile_fpregs_reg_4__0_ ( .D(n7378), .CK(clock), .Q(
        decode_regfile_fpregs_4__0_) );
  DFF_X2 decode_regfile_fpregs_reg_4__1_ ( .D(n7377), .CK(clock), .Q(
        decode_regfile_fpregs_4__1_) );
  DFF_X2 decode_regfile_fpregs_reg_4__2_ ( .D(n7376), .CK(clock), .Q(
        decode_regfile_fpregs_4__2_) );
  DFF_X2 decode_regfile_fpregs_reg_4__3_ ( .D(n7375), .CK(clock), .Q(
        decode_regfile_fpregs_4__3_) );
  DFF_X2 decode_regfile_fpregs_reg_4__4_ ( .D(n7374), .CK(clock), .Q(
        decode_regfile_fpregs_4__4_) );
  DFF_X2 decode_regfile_fpregs_reg_4__5_ ( .D(n7373), .CK(clock), .Q(
        decode_regfile_fpregs_4__5_) );
  DFF_X2 decode_regfile_fpregs_reg_4__6_ ( .D(n7372), .CK(clock), .Q(
        decode_regfile_fpregs_4__6_) );
  DFF_X2 decode_regfile_fpregs_reg_4__7_ ( .D(n7371), .CK(clock), .Q(
        decode_regfile_fpregs_4__7_) );
  DFF_X2 decode_regfile_fpregs_reg_4__8_ ( .D(n7370), .CK(clock), .Q(
        decode_regfile_fpregs_4__8_) );
  DFF_X2 decode_regfile_fpregs_reg_4__9_ ( .D(n7369), .CK(clock), .Q(
        decode_regfile_fpregs_4__9_) );
  DFF_X2 decode_regfile_fpregs_reg_4__10_ ( .D(n7368), .CK(clock), .Q(
        decode_regfile_fpregs_4__10_) );
  DFF_X2 decode_regfile_fpregs_reg_4__11_ ( .D(n7367), .CK(clock), .Q(
        decode_regfile_fpregs_4__11_) );
  DFF_X2 decode_regfile_fpregs_reg_4__12_ ( .D(n7366), .CK(clock), .Q(
        decode_regfile_fpregs_4__12_) );
  DFF_X2 decode_regfile_fpregs_reg_4__13_ ( .D(n7365), .CK(clock), .Q(
        decode_regfile_fpregs_4__13_) );
  DFF_X2 decode_regfile_fpregs_reg_4__14_ ( .D(n7364), .CK(clock), .Q(
        decode_regfile_fpregs_4__14_) );
  DFF_X2 decode_regfile_fpregs_reg_4__15_ ( .D(n7363), .CK(clock), .Q(
        decode_regfile_fpregs_4__15_) );
  DFF_X2 decode_regfile_fpregs_reg_4__16_ ( .D(n7362), .CK(clock), .Q(
        decode_regfile_fpregs_4__16_) );
  DFF_X2 decode_regfile_fpregs_reg_4__17_ ( .D(n7361), .CK(clock), .Q(
        decode_regfile_fpregs_4__17_) );
  DFF_X2 decode_regfile_fpregs_reg_4__18_ ( .D(n7360), .CK(clock), .Q(
        decode_regfile_fpregs_4__18_) );
  DFF_X2 decode_regfile_fpregs_reg_4__19_ ( .D(n7359), .CK(clock), .Q(
        decode_regfile_fpregs_4__19_) );
  DFF_X2 decode_regfile_fpregs_reg_4__20_ ( .D(n7358), .CK(clock), .Q(
        decode_regfile_fpregs_4__20_) );
  DFF_X2 decode_regfile_fpregs_reg_4__21_ ( .D(n7357), .CK(clock), .Q(
        decode_regfile_fpregs_4__21_) );
  DFF_X2 decode_regfile_fpregs_reg_4__22_ ( .D(n7356), .CK(clock), .Q(
        decode_regfile_fpregs_4__22_) );
  DFF_X2 decode_regfile_fpregs_reg_4__23_ ( .D(n7355), .CK(clock), .Q(
        decode_regfile_fpregs_4__23_) );
  DFF_X2 decode_regfile_fpregs_reg_4__24_ ( .D(n7354), .CK(clock), .Q(
        decode_regfile_fpregs_4__24_) );
  DFF_X2 decode_regfile_fpregs_reg_4__25_ ( .D(n7353), .CK(clock), .Q(
        decode_regfile_fpregs_4__25_) );
  DFF_X2 decode_regfile_fpregs_reg_4__26_ ( .D(n7352), .CK(clock), .Q(
        decode_regfile_fpregs_4__26_) );
  DFF_X2 decode_regfile_fpregs_reg_4__27_ ( .D(n7351), .CK(clock), .Q(
        decode_regfile_fpregs_4__27_) );
  DFF_X2 decode_regfile_fpregs_reg_4__28_ ( .D(n7350), .CK(clock), .Q(
        decode_regfile_fpregs_4__28_) );
  DFF_X2 decode_regfile_fpregs_reg_4__29_ ( .D(n7349), .CK(clock), .Q(
        decode_regfile_fpregs_4__29_) );
  DFF_X2 decode_regfile_fpregs_reg_4__30_ ( .D(n7348), .CK(clock), .Q(
        decode_regfile_fpregs_4__30_) );
  DFF_X2 decode_regfile_fpregs_reg_4__31_ ( .D(n7347), .CK(clock), .Q(
        decode_regfile_fpregs_4__31_) );
  DFF_X2 decode_regfile_fpregs_reg_3__0_ ( .D(n7346), .CK(clock), .Q(
        decode_regfile_fpregs_3__0_) );
  DFF_X2 decode_regfile_fpregs_reg_3__1_ ( .D(n7345), .CK(clock), .Q(
        decode_regfile_fpregs_3__1_) );
  DFF_X2 decode_regfile_fpregs_reg_3__2_ ( .D(n7344), .CK(clock), .Q(
        decode_regfile_fpregs_3__2_) );
  DFF_X2 decode_regfile_fpregs_reg_3__3_ ( .D(n7343), .CK(clock), .Q(
        decode_regfile_fpregs_3__3_) );
  DFF_X2 decode_regfile_fpregs_reg_3__4_ ( .D(n7342), .CK(clock), .Q(
        decode_regfile_fpregs_3__4_) );
  DFF_X2 decode_regfile_fpregs_reg_3__5_ ( .D(n7341), .CK(clock), .Q(
        decode_regfile_fpregs_3__5_) );
  DFF_X2 decode_regfile_fpregs_reg_3__6_ ( .D(n7340), .CK(clock), .Q(
        decode_regfile_fpregs_3__6_) );
  DFF_X2 decode_regfile_fpregs_reg_3__7_ ( .D(n7339), .CK(clock), .Q(
        decode_regfile_fpregs_3__7_) );
  DFF_X2 decode_regfile_fpregs_reg_3__8_ ( .D(n7338), .CK(clock), .Q(
        decode_regfile_fpregs_3__8_) );
  DFF_X2 decode_regfile_fpregs_reg_3__9_ ( .D(n7337), .CK(clock), .Q(
        decode_regfile_fpregs_3__9_) );
  DFF_X2 decode_regfile_fpregs_reg_3__10_ ( .D(n7336), .CK(clock), .Q(
        decode_regfile_fpregs_3__10_) );
  DFF_X2 decode_regfile_fpregs_reg_3__11_ ( .D(n7335), .CK(clock), .Q(
        decode_regfile_fpregs_3__11_) );
  DFF_X2 decode_regfile_fpregs_reg_3__12_ ( .D(n7334), .CK(clock), .Q(
        decode_regfile_fpregs_3__12_) );
  DFF_X2 decode_regfile_fpregs_reg_3__13_ ( .D(n7333), .CK(clock), .Q(
        decode_regfile_fpregs_3__13_) );
  DFF_X2 decode_regfile_fpregs_reg_3__14_ ( .D(n7332), .CK(clock), .Q(
        decode_regfile_fpregs_3__14_) );
  DFF_X2 decode_regfile_fpregs_reg_3__15_ ( .D(n7331), .CK(clock), .Q(
        decode_regfile_fpregs_3__15_) );
  DFF_X2 decode_regfile_fpregs_reg_3__16_ ( .D(n7330), .CK(clock), .Q(
        decode_regfile_fpregs_3__16_) );
  DFF_X2 decode_regfile_fpregs_reg_3__17_ ( .D(n7329), .CK(clock), .Q(
        decode_regfile_fpregs_3__17_) );
  DFF_X2 decode_regfile_fpregs_reg_3__18_ ( .D(n7328), .CK(clock), .Q(
        decode_regfile_fpregs_3__18_) );
  DFF_X2 decode_regfile_fpregs_reg_3__19_ ( .D(n7327), .CK(clock), .Q(
        decode_regfile_fpregs_3__19_) );
  DFF_X2 decode_regfile_fpregs_reg_3__20_ ( .D(n7326), .CK(clock), .Q(
        decode_regfile_fpregs_3__20_) );
  DFF_X2 decode_regfile_fpregs_reg_3__21_ ( .D(n7325), .CK(clock), .Q(
        decode_regfile_fpregs_3__21_) );
  DFF_X2 decode_regfile_fpregs_reg_3__22_ ( .D(n7324), .CK(clock), .Q(
        decode_regfile_fpregs_3__22_) );
  DFF_X2 decode_regfile_fpregs_reg_3__23_ ( .D(n7323), .CK(clock), .Q(
        decode_regfile_fpregs_3__23_) );
  DFF_X2 decode_regfile_fpregs_reg_3__24_ ( .D(n7322), .CK(clock), .Q(
        decode_regfile_fpregs_3__24_) );
  DFF_X2 decode_regfile_fpregs_reg_3__25_ ( .D(n7321), .CK(clock), .Q(
        decode_regfile_fpregs_3__25_) );
  DFF_X2 decode_regfile_fpregs_reg_3__26_ ( .D(n7320), .CK(clock), .Q(
        decode_regfile_fpregs_3__26_) );
  DFF_X2 decode_regfile_fpregs_reg_3__27_ ( .D(n7319), .CK(clock), .Q(
        decode_regfile_fpregs_3__27_) );
  DFF_X2 decode_regfile_fpregs_reg_3__28_ ( .D(n7318), .CK(clock), .Q(
        decode_regfile_fpregs_3__28_) );
  DFF_X2 decode_regfile_fpregs_reg_3__29_ ( .D(n7317), .CK(clock), .Q(
        decode_regfile_fpregs_3__29_) );
  DFF_X2 decode_regfile_fpregs_reg_3__30_ ( .D(n7316), .CK(clock), .Q(
        decode_regfile_fpregs_3__30_) );
  DFF_X2 decode_regfile_fpregs_reg_3__31_ ( .D(n7315), .CK(clock), .Q(
        decode_regfile_fpregs_3__31_) );
  DFF_X2 decode_regfile_fpregs_reg_2__0_ ( .D(n7314), .CK(clock), .Q(
        decode_regfile_fpregs_2__0_) );
  DFF_X2 decode_regfile_fpregs_reg_2__1_ ( .D(n7313), .CK(clock), .Q(
        decode_regfile_fpregs_2__1_) );
  DFF_X2 decode_regfile_fpregs_reg_2__2_ ( .D(n7312), .CK(clock), .Q(
        decode_regfile_fpregs_2__2_) );
  DFF_X2 decode_regfile_fpregs_reg_2__3_ ( .D(n7311), .CK(clock), .Q(
        decode_regfile_fpregs_2__3_) );
  DFF_X2 decode_regfile_fpregs_reg_2__4_ ( .D(n7310), .CK(clock), .Q(
        decode_regfile_fpregs_2__4_) );
  DFF_X2 decode_regfile_fpregs_reg_2__5_ ( .D(n7309), .CK(clock), .Q(
        decode_regfile_fpregs_2__5_) );
  DFF_X2 decode_regfile_fpregs_reg_2__6_ ( .D(n7308), .CK(clock), .Q(
        decode_regfile_fpregs_2__6_) );
  DFF_X2 decode_regfile_fpregs_reg_2__7_ ( .D(n7307), .CK(clock), .Q(
        decode_regfile_fpregs_2__7_) );
  DFF_X2 decode_regfile_fpregs_reg_2__8_ ( .D(n7306), .CK(clock), .Q(
        decode_regfile_fpregs_2__8_) );
  DFF_X2 decode_regfile_fpregs_reg_2__9_ ( .D(n7305), .CK(clock), .Q(
        decode_regfile_fpregs_2__9_) );
  DFF_X2 decode_regfile_fpregs_reg_2__10_ ( .D(n7304), .CK(clock), .Q(
        decode_regfile_fpregs_2__10_) );
  DFF_X2 decode_regfile_fpregs_reg_2__11_ ( .D(n7303), .CK(clock), .Q(
        decode_regfile_fpregs_2__11_) );
  DFF_X2 decode_regfile_fpregs_reg_2__12_ ( .D(n7302), .CK(clock), .Q(
        decode_regfile_fpregs_2__12_) );
  DFF_X2 decode_regfile_fpregs_reg_2__13_ ( .D(n7301), .CK(clock), .Q(
        decode_regfile_fpregs_2__13_) );
  DFF_X2 decode_regfile_fpregs_reg_2__14_ ( .D(n7300), .CK(clock), .Q(
        decode_regfile_fpregs_2__14_) );
  DFF_X2 decode_regfile_fpregs_reg_2__15_ ( .D(n7299), .CK(clock), .Q(
        decode_regfile_fpregs_2__15_) );
  DFF_X2 decode_regfile_fpregs_reg_2__16_ ( .D(n7298), .CK(clock), .Q(
        decode_regfile_fpregs_2__16_) );
  DFF_X2 decode_regfile_fpregs_reg_2__17_ ( .D(n7297), .CK(clock), .Q(
        decode_regfile_fpregs_2__17_) );
  DFF_X2 decode_regfile_fpregs_reg_2__18_ ( .D(n7296), .CK(clock), .Q(
        decode_regfile_fpregs_2__18_) );
  DFF_X2 decode_regfile_fpregs_reg_2__19_ ( .D(n7295), .CK(clock), .Q(
        decode_regfile_fpregs_2__19_) );
  DFF_X2 decode_regfile_fpregs_reg_2__20_ ( .D(n7294), .CK(clock), .Q(
        decode_regfile_fpregs_2__20_) );
  DFF_X2 decode_regfile_fpregs_reg_2__21_ ( .D(n7293), .CK(clock), .Q(
        decode_regfile_fpregs_2__21_) );
  DFF_X2 decode_regfile_fpregs_reg_2__22_ ( .D(n7292), .CK(clock), .Q(
        decode_regfile_fpregs_2__22_) );
  DFF_X2 decode_regfile_fpregs_reg_2__23_ ( .D(n7291), .CK(clock), .Q(
        decode_regfile_fpregs_2__23_) );
  DFF_X2 decode_regfile_fpregs_reg_2__24_ ( .D(n7290), .CK(clock), .Q(
        decode_regfile_fpregs_2__24_) );
  DFF_X2 decode_regfile_fpregs_reg_2__25_ ( .D(n7289), .CK(clock), .Q(
        decode_regfile_fpregs_2__25_) );
  DFF_X2 decode_regfile_fpregs_reg_2__26_ ( .D(n7288), .CK(clock), .Q(
        decode_regfile_fpregs_2__26_) );
  DFF_X2 decode_regfile_fpregs_reg_2__27_ ( .D(n7287), .CK(clock), .Q(
        decode_regfile_fpregs_2__27_) );
  DFF_X2 decode_regfile_fpregs_reg_2__28_ ( .D(n7286), .CK(clock), .Q(
        decode_regfile_fpregs_2__28_) );
  DFF_X2 decode_regfile_fpregs_reg_2__29_ ( .D(n7285), .CK(clock), .Q(
        decode_regfile_fpregs_2__29_) );
  DFF_X2 decode_regfile_fpregs_reg_2__30_ ( .D(n7284), .CK(clock), .Q(
        decode_regfile_fpregs_2__30_) );
  DFF_X2 decode_regfile_fpregs_reg_2__31_ ( .D(n7283), .CK(clock), .Q(
        decode_regfile_fpregs_2__31_) );
  DFF_X2 decode_regfile_fpregs_reg_1__0_ ( .D(n7282), .CK(clock), .Q(
        decode_regfile_fpregs_1__0_) );
  DFF_X2 decode_regfile_fpregs_reg_1__1_ ( .D(n7281), .CK(clock), .Q(
        decode_regfile_fpregs_1__1_) );
  DFF_X2 decode_regfile_fpregs_reg_1__2_ ( .D(n7280), .CK(clock), .Q(
        decode_regfile_fpregs_1__2_) );
  DFF_X2 decode_regfile_fpregs_reg_1__3_ ( .D(n7279), .CK(clock), .Q(
        decode_regfile_fpregs_1__3_) );
  DFF_X2 decode_regfile_fpregs_reg_1__4_ ( .D(n7278), .CK(clock), .Q(
        decode_regfile_fpregs_1__4_) );
  DFF_X2 decode_regfile_fpregs_reg_1__5_ ( .D(n7277), .CK(clock), .Q(
        decode_regfile_fpregs_1__5_) );
  DFF_X2 decode_regfile_fpregs_reg_1__6_ ( .D(n7276), .CK(clock), .Q(
        decode_regfile_fpregs_1__6_) );
  DFF_X2 decode_regfile_fpregs_reg_1__7_ ( .D(n7275), .CK(clock), .Q(
        decode_regfile_fpregs_1__7_) );
  DFF_X2 decode_regfile_fpregs_reg_1__8_ ( .D(n7274), .CK(clock), .Q(
        decode_regfile_fpregs_1__8_) );
  DFF_X2 decode_regfile_fpregs_reg_1__9_ ( .D(n7273), .CK(clock), .Q(
        decode_regfile_fpregs_1__9_) );
  DFF_X2 decode_regfile_fpregs_reg_1__10_ ( .D(n7272), .CK(clock), .Q(
        decode_regfile_fpregs_1__10_) );
  DFF_X2 decode_regfile_fpregs_reg_1__11_ ( .D(n7271), .CK(clock), .Q(
        decode_regfile_fpregs_1__11_) );
  DFF_X2 decode_regfile_fpregs_reg_1__12_ ( .D(n7270), .CK(clock), .Q(
        decode_regfile_fpregs_1__12_) );
  DFF_X2 decode_regfile_fpregs_reg_1__13_ ( .D(n7269), .CK(clock), .Q(
        decode_regfile_fpregs_1__13_) );
  DFF_X2 decode_regfile_fpregs_reg_1__14_ ( .D(n7268), .CK(clock), .Q(
        decode_regfile_fpregs_1__14_) );
  DFF_X2 decode_regfile_fpregs_reg_1__15_ ( .D(n7267), .CK(clock), .Q(
        decode_regfile_fpregs_1__15_) );
  DFF_X2 decode_regfile_fpregs_reg_1__16_ ( .D(n7266), .CK(clock), .Q(
        decode_regfile_fpregs_1__16_) );
  DFF_X2 decode_regfile_fpregs_reg_1__17_ ( .D(n7265), .CK(clock), .Q(
        decode_regfile_fpregs_1__17_) );
  DFF_X2 decode_regfile_fpregs_reg_1__18_ ( .D(n7264), .CK(clock), .Q(
        decode_regfile_fpregs_1__18_) );
  DFF_X2 decode_regfile_fpregs_reg_1__19_ ( .D(n7263), .CK(clock), .Q(
        decode_regfile_fpregs_1__19_) );
  DFF_X2 decode_regfile_fpregs_reg_1__20_ ( .D(n7262), .CK(clock), .Q(
        decode_regfile_fpregs_1__20_) );
  DFF_X2 decode_regfile_fpregs_reg_1__21_ ( .D(n7261), .CK(clock), .Q(
        decode_regfile_fpregs_1__21_) );
  DFF_X2 decode_regfile_fpregs_reg_1__22_ ( .D(n7260), .CK(clock), .Q(
        decode_regfile_fpregs_1__22_) );
  DFF_X2 decode_regfile_fpregs_reg_1__23_ ( .D(n7259), .CK(clock), .Q(
        decode_regfile_fpregs_1__23_) );
  DFF_X2 decode_regfile_fpregs_reg_1__24_ ( .D(n7258), .CK(clock), .Q(
        decode_regfile_fpregs_1__24_) );
  DFF_X2 decode_regfile_fpregs_reg_1__25_ ( .D(n7257), .CK(clock), .Q(
        decode_regfile_fpregs_1__25_) );
  DFF_X2 decode_regfile_fpregs_reg_1__26_ ( .D(n7256), .CK(clock), .Q(
        decode_regfile_fpregs_1__26_) );
  DFF_X2 decode_regfile_fpregs_reg_1__27_ ( .D(n7255), .CK(clock), .Q(
        decode_regfile_fpregs_1__27_) );
  DFF_X2 decode_regfile_fpregs_reg_1__28_ ( .D(n7254), .CK(clock), .Q(
        decode_regfile_fpregs_1__28_) );
  DFF_X2 decode_regfile_fpregs_reg_1__29_ ( .D(n7253), .CK(clock), .Q(
        decode_regfile_fpregs_1__29_) );
  DFF_X2 decode_regfile_fpregs_reg_1__30_ ( .D(n7252), .CK(clock), .Q(
        decode_regfile_fpregs_1__30_) );
  DFF_X2 decode_regfile_fpregs_reg_1__31_ ( .D(n7251), .CK(clock), .Q(
        decode_regfile_fpregs_1__31_) );
  DFF_X2 decode_regfile_fpregs_reg_0__0_ ( .D(n7250), .CK(clock), .Q(
        decode_regfile_fpregs_0__0_) );
  DFF_X2 decode_regfile_fpregs_reg_0__1_ ( .D(n7249), .CK(clock), .Q(
        decode_regfile_fpregs_0__1_) );
  DFF_X2 decode_regfile_fpregs_reg_0__2_ ( .D(n7248), .CK(clock), .Q(
        decode_regfile_fpregs_0__2_) );
  DFF_X2 decode_regfile_fpregs_reg_0__3_ ( .D(n7247), .CK(clock), .Q(
        decode_regfile_fpregs_0__3_) );
  DFF_X2 decode_regfile_fpregs_reg_0__4_ ( .D(n7246), .CK(clock), .Q(
        decode_regfile_fpregs_0__4_) );
  DFF_X2 decode_regfile_fpregs_reg_0__5_ ( .D(n7245), .CK(clock), .Q(
        decode_regfile_fpregs_0__5_) );
  DFF_X2 decode_regfile_fpregs_reg_0__6_ ( .D(n7244), .CK(clock), .Q(
        decode_regfile_fpregs_0__6_) );
  DFF_X2 decode_regfile_fpregs_reg_0__7_ ( .D(n7243), .CK(clock), .Q(
        decode_regfile_fpregs_0__7_) );
  DFF_X2 decode_regfile_fpregs_reg_0__8_ ( .D(n7242), .CK(clock), .Q(
        decode_regfile_fpregs_0__8_) );
  DFF_X2 decode_regfile_fpregs_reg_0__9_ ( .D(n7241), .CK(clock), .Q(
        decode_regfile_fpregs_0__9_) );
  DFF_X2 decode_regfile_fpregs_reg_0__10_ ( .D(n7240), .CK(clock), .Q(
        decode_regfile_fpregs_0__10_) );
  DFF_X2 decode_regfile_fpregs_reg_0__11_ ( .D(n7239), .CK(clock), .Q(
        decode_regfile_fpregs_0__11_) );
  DFF_X2 decode_regfile_fpregs_reg_0__12_ ( .D(n7238), .CK(clock), .Q(
        decode_regfile_fpregs_0__12_) );
  DFF_X2 decode_regfile_fpregs_reg_0__13_ ( .D(n7237), .CK(clock), .Q(
        decode_regfile_fpregs_0__13_) );
  DFF_X2 decode_regfile_fpregs_reg_0__14_ ( .D(n7236), .CK(clock), .Q(
        decode_regfile_fpregs_0__14_) );
  DFF_X2 decode_regfile_fpregs_reg_0__15_ ( .D(n7235), .CK(clock), .Q(
        decode_regfile_fpregs_0__15_) );
  DFF_X2 decode_regfile_fpregs_reg_0__16_ ( .D(n7234), .CK(clock), .Q(
        decode_regfile_fpregs_0__16_) );
  DFF_X2 decode_regfile_fpregs_reg_0__17_ ( .D(n7233), .CK(clock), .Q(
        decode_regfile_fpregs_0__17_) );
  DFF_X2 decode_regfile_fpregs_reg_0__18_ ( .D(n7232), .CK(clock), .Q(
        decode_regfile_fpregs_0__18_) );
  DFF_X2 decode_regfile_fpregs_reg_0__19_ ( .D(n7231), .CK(clock), .Q(
        decode_regfile_fpregs_0__19_) );
  DFF_X2 decode_regfile_fpregs_reg_0__20_ ( .D(n7230), .CK(clock), .Q(
        decode_regfile_fpregs_0__20_) );
  DFF_X2 decode_regfile_fpregs_reg_0__21_ ( .D(n7229), .CK(clock), .Q(
        decode_regfile_fpregs_0__21_) );
  DFF_X2 decode_regfile_fpregs_reg_0__22_ ( .D(n7228), .CK(clock), .Q(
        decode_regfile_fpregs_0__22_) );
  DFF_X2 decode_regfile_fpregs_reg_0__23_ ( .D(n7227), .CK(clock), .Q(
        decode_regfile_fpregs_0__23_) );
  DFF_X2 decode_regfile_fpregs_reg_0__24_ ( .D(n7226), .CK(clock), .Q(
        decode_regfile_fpregs_0__24_) );
  DFF_X2 decode_regfile_fpregs_reg_0__25_ ( .D(n7225), .CK(clock), .Q(
        decode_regfile_fpregs_0__25_) );
  DFF_X2 decode_regfile_fpregs_reg_0__26_ ( .D(n7224), .CK(clock), .Q(
        decode_regfile_fpregs_0__26_) );
  DFF_X2 decode_regfile_fpregs_reg_0__27_ ( .D(n7223), .CK(clock), .Q(
        decode_regfile_fpregs_0__27_) );
  DFF_X2 decode_regfile_fpregs_reg_0__28_ ( .D(n7222), .CK(clock), .Q(
        decode_regfile_fpregs_0__28_) );
  DFF_X2 decode_regfile_fpregs_reg_0__29_ ( .D(n7221), .CK(clock), .Q(
        decode_regfile_fpregs_0__29_) );
  DFF_X2 decode_regfile_fpregs_reg_0__30_ ( .D(n7220), .CK(clock), .Q(
        decode_regfile_fpregs_0__30_) );
  DFF_X2 decode_regfile_fpregs_reg_0__31_ ( .D(n7219), .CK(clock), .Q(
        decode_regfile_fpregs_0__31_) );
  DFF_X2 decode_regfile_intregs_reg_31__0_ ( .D(n7218), .CK(clock), .Q(
        decode_regfile_intregs_31__0_) );
  DFF_X2 decode_regfile_intregs_reg_31__1_ ( .D(n7217), .CK(clock), .Q(
        decode_regfile_intregs_31__1_) );
  DFF_X2 decode_regfile_intregs_reg_31__2_ ( .D(n7216), .CK(clock), .Q(
        decode_regfile_intregs_31__2_) );
  DFF_X2 decode_regfile_intregs_reg_31__3_ ( .D(n7215), .CK(clock), .Q(
        decode_regfile_intregs_31__3_) );
  DFF_X2 decode_regfile_intregs_reg_31__4_ ( .D(n7214), .CK(clock), .Q(
        decode_regfile_intregs_31__4_) );
  DFF_X2 decode_regfile_intregs_reg_31__5_ ( .D(n7213), .CK(clock), .Q(
        decode_regfile_intregs_31__5_) );
  DFF_X2 decode_regfile_intregs_reg_31__6_ ( .D(n7212), .CK(clock), .Q(
        decode_regfile_intregs_31__6_) );
  DFF_X2 decode_regfile_intregs_reg_31__7_ ( .D(n7211), .CK(clock), .Q(
        decode_regfile_intregs_31__7_) );
  DFF_X2 decode_regfile_intregs_reg_31__8_ ( .D(n7210), .CK(clock), .Q(
        decode_regfile_intregs_31__8_) );
  DFF_X2 decode_regfile_intregs_reg_31__9_ ( .D(n7209), .CK(clock), .Q(
        decode_regfile_intregs_31__9_) );
  DFF_X2 decode_regfile_intregs_reg_31__10_ ( .D(n7208), .CK(clock), .Q(
        decode_regfile_intregs_31__10_) );
  DFF_X2 decode_regfile_intregs_reg_31__11_ ( .D(n7207), .CK(clock), .Q(
        decode_regfile_intregs_31__11_) );
  DFF_X2 decode_regfile_intregs_reg_31__12_ ( .D(n7206), .CK(clock), .Q(
        decode_regfile_intregs_31__12_) );
  DFF_X2 decode_regfile_intregs_reg_31__13_ ( .D(n7205), .CK(clock), .Q(
        decode_regfile_intregs_31__13_) );
  DFF_X2 decode_regfile_intregs_reg_31__14_ ( .D(n7204), .CK(clock), .Q(
        decode_regfile_intregs_31__14_) );
  DFF_X2 decode_regfile_intregs_reg_31__15_ ( .D(n7203), .CK(clock), .Q(
        decode_regfile_intregs_31__15_) );
  DFF_X2 decode_regfile_intregs_reg_31__16_ ( .D(n7202), .CK(clock), .Q(
        decode_regfile_intregs_31__16_) );
  DFF_X2 decode_regfile_intregs_reg_31__17_ ( .D(n7201), .CK(clock), .Q(
        decode_regfile_intregs_31__17_) );
  DFF_X2 decode_regfile_intregs_reg_31__18_ ( .D(n7200), .CK(clock), .Q(
        decode_regfile_intregs_31__18_) );
  DFF_X2 decode_regfile_intregs_reg_31__19_ ( .D(n7199), .CK(clock), .Q(
        decode_regfile_intregs_31__19_) );
  DFF_X2 decode_regfile_intregs_reg_31__20_ ( .D(n7198), .CK(clock), .Q(
        decode_regfile_intregs_31__20_) );
  DFF_X2 decode_regfile_intregs_reg_31__21_ ( .D(n7197), .CK(clock), .Q(
        decode_regfile_intregs_31__21_) );
  DFF_X2 decode_regfile_intregs_reg_31__22_ ( .D(n7196), .CK(clock), .Q(
        decode_regfile_intregs_31__22_) );
  DFF_X2 decode_regfile_intregs_reg_31__23_ ( .D(n7195), .CK(clock), .Q(
        decode_regfile_intregs_31__23_) );
  DFF_X2 decode_regfile_intregs_reg_31__24_ ( .D(n7194), .CK(clock), .Q(
        decode_regfile_intregs_31__24_) );
  DFF_X2 decode_regfile_intregs_reg_31__25_ ( .D(n7193), .CK(clock), .Q(
        decode_regfile_intregs_31__25_) );
  DFF_X2 decode_regfile_intregs_reg_31__26_ ( .D(n7192), .CK(clock), .Q(
        decode_regfile_intregs_31__26_) );
  DFF_X2 decode_regfile_intregs_reg_31__27_ ( .D(n7191), .CK(clock), .Q(
        decode_regfile_intregs_31__27_) );
  DFF_X2 decode_regfile_intregs_reg_31__28_ ( .D(n7190), .CK(clock), .Q(
        decode_regfile_intregs_31__28_) );
  DFF_X2 decode_regfile_intregs_reg_31__29_ ( .D(n7189), .CK(clock), .Q(
        decode_regfile_intregs_31__29_) );
  DFF_X2 decode_regfile_intregs_reg_31__30_ ( .D(n7188), .CK(clock), .Q(
        decode_regfile_intregs_31__30_) );
  DFF_X2 decode_regfile_intregs_reg_31__31_ ( .D(n7187), .CK(clock), .Q(
        decode_regfile_intregs_31__31_) );
  DFF_X2 decode_regfile_intregs_reg_30__0_ ( .D(n7186), .CK(clock), .Q(
        decode_regfile_intregs_30__0_) );
  DFF_X2 decode_regfile_intregs_reg_30__1_ ( .D(n7185), .CK(clock), .Q(
        decode_regfile_intregs_30__1_) );
  DFF_X2 decode_regfile_intregs_reg_30__2_ ( .D(n7184), .CK(clock), .Q(
        decode_regfile_intregs_30__2_) );
  DFF_X2 decode_regfile_intregs_reg_30__3_ ( .D(n7183), .CK(clock), .Q(
        decode_regfile_intregs_30__3_) );
  DFF_X2 decode_regfile_intregs_reg_30__4_ ( .D(n7182), .CK(clock), .Q(
        decode_regfile_intregs_30__4_) );
  DFF_X2 decode_regfile_intregs_reg_30__5_ ( .D(n7181), .CK(clock), .Q(
        decode_regfile_intregs_30__5_) );
  DFF_X2 decode_regfile_intregs_reg_30__6_ ( .D(n7180), .CK(clock), .Q(
        decode_regfile_intregs_30__6_) );
  DFF_X2 decode_regfile_intregs_reg_30__7_ ( .D(n7179), .CK(clock), .Q(
        decode_regfile_intregs_30__7_) );
  DFF_X2 decode_regfile_intregs_reg_30__8_ ( .D(n7178), .CK(clock), .Q(
        decode_regfile_intregs_30__8_) );
  DFF_X2 decode_regfile_intregs_reg_30__9_ ( .D(n7177), .CK(clock), .Q(
        decode_regfile_intregs_30__9_) );
  DFF_X2 decode_regfile_intregs_reg_30__10_ ( .D(n7176), .CK(clock), .Q(
        decode_regfile_intregs_30__10_) );
  DFF_X2 decode_regfile_intregs_reg_30__11_ ( .D(n7175), .CK(clock), .Q(
        decode_regfile_intregs_30__11_) );
  DFF_X2 decode_regfile_intregs_reg_30__12_ ( .D(n7174), .CK(clock), .Q(
        decode_regfile_intregs_30__12_) );
  DFF_X2 decode_regfile_intregs_reg_30__13_ ( .D(n7173), .CK(clock), .Q(
        decode_regfile_intregs_30__13_) );
  DFF_X2 decode_regfile_intregs_reg_30__14_ ( .D(n7172), .CK(clock), .Q(
        decode_regfile_intregs_30__14_) );
  DFF_X2 decode_regfile_intregs_reg_30__15_ ( .D(n7171), .CK(clock), .Q(
        decode_regfile_intregs_30__15_) );
  DFF_X2 decode_regfile_intregs_reg_30__16_ ( .D(n7170), .CK(clock), .Q(
        decode_regfile_intregs_30__16_) );
  DFF_X2 decode_regfile_intregs_reg_30__17_ ( .D(n7169), .CK(clock), .Q(
        decode_regfile_intregs_30__17_) );
  DFF_X2 decode_regfile_intregs_reg_30__18_ ( .D(n7168), .CK(clock), .Q(
        decode_regfile_intregs_30__18_) );
  DFF_X2 decode_regfile_intregs_reg_30__19_ ( .D(n7167), .CK(clock), .Q(
        decode_regfile_intregs_30__19_) );
  DFF_X2 decode_regfile_intregs_reg_30__20_ ( .D(n7166), .CK(clock), .Q(
        decode_regfile_intregs_30__20_) );
  DFF_X2 decode_regfile_intregs_reg_30__21_ ( .D(n7165), .CK(clock), .Q(
        decode_regfile_intregs_30__21_) );
  DFF_X2 decode_regfile_intregs_reg_30__22_ ( .D(n7164), .CK(clock), .Q(
        decode_regfile_intregs_30__22_) );
  DFF_X2 decode_regfile_intregs_reg_30__23_ ( .D(n7163), .CK(clock), .Q(
        decode_regfile_intregs_30__23_) );
  DFF_X2 decode_regfile_intregs_reg_30__24_ ( .D(n7162), .CK(clock), .Q(
        decode_regfile_intregs_30__24_) );
  DFF_X2 decode_regfile_intregs_reg_30__25_ ( .D(n7161), .CK(clock), .Q(
        decode_regfile_intregs_30__25_) );
  DFF_X2 decode_regfile_intregs_reg_30__26_ ( .D(n7160), .CK(clock), .Q(
        decode_regfile_intregs_30__26_) );
  DFF_X2 decode_regfile_intregs_reg_30__27_ ( .D(n7159), .CK(clock), .Q(
        decode_regfile_intregs_30__27_) );
  DFF_X2 decode_regfile_intregs_reg_30__28_ ( .D(n7158), .CK(clock), .Q(
        decode_regfile_intregs_30__28_) );
  DFF_X2 decode_regfile_intregs_reg_30__29_ ( .D(n7157), .CK(clock), .Q(
        decode_regfile_intregs_30__29_) );
  DFF_X2 decode_regfile_intregs_reg_30__30_ ( .D(n7156), .CK(clock), .Q(
        decode_regfile_intregs_30__30_) );
  DFF_X2 decode_regfile_intregs_reg_30__31_ ( .D(n7155), .CK(clock), .Q(
        decode_regfile_intregs_30__31_) );
  DFF_X2 decode_regfile_intregs_reg_29__0_ ( .D(n7154), .CK(clock), .Q(
        decode_regfile_intregs_29__0_) );
  DFF_X2 decode_regfile_intregs_reg_29__1_ ( .D(n7153), .CK(clock), .Q(
        decode_regfile_intregs_29__1_) );
  DFF_X2 decode_regfile_intregs_reg_29__2_ ( .D(n7152), .CK(clock), .Q(
        decode_regfile_intregs_29__2_) );
  DFF_X2 decode_regfile_intregs_reg_29__3_ ( .D(n7151), .CK(clock), .Q(
        decode_regfile_intregs_29__3_) );
  DFF_X2 decode_regfile_intregs_reg_29__4_ ( .D(n7150), .CK(clock), .Q(
        decode_regfile_intregs_29__4_) );
  DFF_X2 decode_regfile_intregs_reg_29__5_ ( .D(n7149), .CK(clock), .Q(
        decode_regfile_intregs_29__5_) );
  DFF_X2 decode_regfile_intregs_reg_29__6_ ( .D(n7148), .CK(clock), .Q(
        decode_regfile_intregs_29__6_) );
  DFF_X2 decode_regfile_intregs_reg_29__7_ ( .D(n7147), .CK(clock), .Q(
        decode_regfile_intregs_29__7_) );
  DFF_X2 decode_regfile_intregs_reg_29__8_ ( .D(n7146), .CK(clock), .Q(
        decode_regfile_intregs_29__8_) );
  DFF_X2 decode_regfile_intregs_reg_29__9_ ( .D(n7145), .CK(clock), .Q(
        decode_regfile_intregs_29__9_) );
  DFF_X2 decode_regfile_intregs_reg_29__10_ ( .D(n7144), .CK(clock), .Q(
        decode_regfile_intregs_29__10_) );
  DFF_X2 decode_regfile_intregs_reg_29__11_ ( .D(n7143), .CK(clock), .Q(
        decode_regfile_intregs_29__11_) );
  DFF_X2 decode_regfile_intregs_reg_29__12_ ( .D(n7142), .CK(clock), .Q(
        decode_regfile_intregs_29__12_) );
  DFF_X2 decode_regfile_intregs_reg_29__13_ ( .D(n7141), .CK(clock), .Q(
        decode_regfile_intregs_29__13_) );
  DFF_X2 decode_regfile_intregs_reg_29__14_ ( .D(n7140), .CK(clock), .Q(
        decode_regfile_intregs_29__14_) );
  DFF_X2 decode_regfile_intregs_reg_29__15_ ( .D(n7139), .CK(clock), .Q(
        decode_regfile_intregs_29__15_) );
  DFF_X2 decode_regfile_intregs_reg_29__16_ ( .D(n7138), .CK(clock), .Q(
        decode_regfile_intregs_29__16_) );
  DFF_X2 decode_regfile_intregs_reg_29__17_ ( .D(n7137), .CK(clock), .Q(
        decode_regfile_intregs_29__17_) );
  DFF_X2 decode_regfile_intregs_reg_29__18_ ( .D(n7136), .CK(clock), .Q(
        decode_regfile_intregs_29__18_) );
  DFF_X2 decode_regfile_intregs_reg_29__19_ ( .D(n7135), .CK(clock), .Q(
        decode_regfile_intregs_29__19_) );
  DFF_X2 decode_regfile_intregs_reg_29__20_ ( .D(n7134), .CK(clock), .Q(
        decode_regfile_intregs_29__20_) );
  DFF_X2 decode_regfile_intregs_reg_29__21_ ( .D(n7133), .CK(clock), .Q(
        decode_regfile_intregs_29__21_) );
  DFF_X2 decode_regfile_intregs_reg_29__22_ ( .D(n7132), .CK(clock), .Q(
        decode_regfile_intregs_29__22_) );
  DFF_X2 decode_regfile_intregs_reg_29__23_ ( .D(n7131), .CK(clock), .Q(
        decode_regfile_intregs_29__23_) );
  DFF_X2 decode_regfile_intregs_reg_29__24_ ( .D(n7130), .CK(clock), .Q(
        decode_regfile_intregs_29__24_) );
  DFF_X2 decode_regfile_intregs_reg_29__25_ ( .D(n7129), .CK(clock), .Q(
        decode_regfile_intregs_29__25_) );
  DFF_X2 decode_regfile_intregs_reg_29__26_ ( .D(n7128), .CK(clock), .Q(
        decode_regfile_intregs_29__26_) );
  DFF_X2 decode_regfile_intregs_reg_29__27_ ( .D(n7127), .CK(clock), .Q(
        decode_regfile_intregs_29__27_) );
  DFF_X2 decode_regfile_intregs_reg_29__28_ ( .D(n7126), .CK(clock), .Q(
        decode_regfile_intregs_29__28_) );
  DFF_X2 decode_regfile_intregs_reg_29__29_ ( .D(n7125), .CK(clock), .Q(
        decode_regfile_intregs_29__29_) );
  DFF_X2 decode_regfile_intregs_reg_29__30_ ( .D(n7124), .CK(clock), .Q(
        decode_regfile_intregs_29__30_) );
  DFF_X2 decode_regfile_intregs_reg_29__31_ ( .D(n7123), .CK(clock), .Q(
        decode_regfile_intregs_29__31_) );
  DFF_X2 decode_regfile_intregs_reg_28__0_ ( .D(n7122), .CK(clock), .Q(
        decode_regfile_intregs_28__0_) );
  DFF_X2 decode_regfile_intregs_reg_28__1_ ( .D(n7121), .CK(clock), .Q(
        decode_regfile_intregs_28__1_) );
  DFF_X2 decode_regfile_intregs_reg_28__2_ ( .D(n7120), .CK(clock), .Q(
        decode_regfile_intregs_28__2_) );
  DFF_X2 decode_regfile_intregs_reg_28__3_ ( .D(n7119), .CK(clock), .Q(
        decode_regfile_intregs_28__3_) );
  DFF_X2 decode_regfile_intregs_reg_28__4_ ( .D(n7118), .CK(clock), .Q(
        decode_regfile_intregs_28__4_) );
  DFF_X2 decode_regfile_intregs_reg_28__5_ ( .D(n7117), .CK(clock), .Q(
        decode_regfile_intregs_28__5_) );
  DFF_X2 decode_regfile_intregs_reg_28__6_ ( .D(n7116), .CK(clock), .Q(
        decode_regfile_intregs_28__6_) );
  DFF_X2 decode_regfile_intregs_reg_28__7_ ( .D(n7115), .CK(clock), .Q(
        decode_regfile_intregs_28__7_) );
  DFF_X2 decode_regfile_intregs_reg_28__8_ ( .D(n7114), .CK(clock), .Q(
        decode_regfile_intregs_28__8_) );
  DFF_X2 decode_regfile_intregs_reg_28__9_ ( .D(n7113), .CK(clock), .Q(
        decode_regfile_intregs_28__9_) );
  DFF_X2 decode_regfile_intregs_reg_28__10_ ( .D(n7112), .CK(clock), .Q(
        decode_regfile_intregs_28__10_) );
  DFF_X2 decode_regfile_intregs_reg_28__11_ ( .D(n7111), .CK(clock), .Q(
        decode_regfile_intregs_28__11_) );
  DFF_X2 decode_regfile_intregs_reg_28__12_ ( .D(n7110), .CK(clock), .Q(
        decode_regfile_intregs_28__12_) );
  DFF_X2 decode_regfile_intregs_reg_28__13_ ( .D(n7109), .CK(clock), .Q(
        decode_regfile_intregs_28__13_) );
  DFF_X2 decode_regfile_intregs_reg_28__14_ ( .D(n7108), .CK(clock), .Q(
        decode_regfile_intregs_28__14_) );
  DFF_X2 decode_regfile_intregs_reg_28__15_ ( .D(n7107), .CK(clock), .Q(
        decode_regfile_intregs_28__15_) );
  DFF_X2 decode_regfile_intregs_reg_28__16_ ( .D(n7106), .CK(clock), .Q(
        decode_regfile_intregs_28__16_) );
  DFF_X2 decode_regfile_intregs_reg_28__17_ ( .D(n7105), .CK(clock), .Q(
        decode_regfile_intregs_28__17_) );
  DFF_X2 decode_regfile_intregs_reg_28__18_ ( .D(n7104), .CK(clock), .Q(
        decode_regfile_intregs_28__18_) );
  DFF_X2 decode_regfile_intregs_reg_28__19_ ( .D(n7103), .CK(clock), .Q(
        decode_regfile_intregs_28__19_) );
  DFF_X2 decode_regfile_intregs_reg_28__20_ ( .D(n7102), .CK(clock), .Q(
        decode_regfile_intregs_28__20_) );
  DFF_X2 decode_regfile_intregs_reg_28__21_ ( .D(n7101), .CK(clock), .Q(
        decode_regfile_intregs_28__21_) );
  DFF_X2 decode_regfile_intregs_reg_28__22_ ( .D(n7100), .CK(clock), .Q(
        decode_regfile_intregs_28__22_) );
  DFF_X2 decode_regfile_intregs_reg_28__23_ ( .D(n7099), .CK(clock), .Q(
        decode_regfile_intregs_28__23_) );
  DFF_X2 decode_regfile_intregs_reg_28__24_ ( .D(n7098), .CK(clock), .Q(
        decode_regfile_intregs_28__24_) );
  DFF_X2 decode_regfile_intregs_reg_28__25_ ( .D(n7097), .CK(clock), .Q(
        decode_regfile_intregs_28__25_) );
  DFF_X2 decode_regfile_intregs_reg_28__26_ ( .D(n7096), .CK(clock), .Q(
        decode_regfile_intregs_28__26_) );
  DFF_X2 decode_regfile_intregs_reg_28__27_ ( .D(n7095), .CK(clock), .Q(
        decode_regfile_intregs_28__27_) );
  DFF_X2 decode_regfile_intregs_reg_28__28_ ( .D(n7094), .CK(clock), .Q(
        decode_regfile_intregs_28__28_) );
  DFF_X2 decode_regfile_intregs_reg_28__29_ ( .D(n7093), .CK(clock), .Q(
        decode_regfile_intregs_28__29_) );
  DFF_X2 decode_regfile_intregs_reg_28__30_ ( .D(n7092), .CK(clock), .Q(
        decode_regfile_intregs_28__30_) );
  DFF_X2 decode_regfile_intregs_reg_28__31_ ( .D(n7091), .CK(clock), .Q(
        decode_regfile_intregs_28__31_) );
  DFF_X2 decode_regfile_intregs_reg_27__0_ ( .D(n7090), .CK(clock), .Q(
        decode_regfile_intregs_27__0_) );
  DFF_X2 decode_regfile_intregs_reg_27__1_ ( .D(n7089), .CK(clock), .Q(
        decode_regfile_intregs_27__1_) );
  DFF_X2 decode_regfile_intregs_reg_27__2_ ( .D(n7088), .CK(clock), .Q(
        decode_regfile_intregs_27__2_) );
  DFF_X2 decode_regfile_intregs_reg_27__3_ ( .D(n7087), .CK(clock), .Q(
        decode_regfile_intregs_27__3_) );
  DFF_X2 decode_regfile_intregs_reg_27__4_ ( .D(n7086), .CK(clock), .Q(
        decode_regfile_intregs_27__4_) );
  DFF_X2 decode_regfile_intregs_reg_27__5_ ( .D(n7085), .CK(clock), .Q(
        decode_regfile_intregs_27__5_) );
  DFF_X2 decode_regfile_intregs_reg_27__6_ ( .D(n7084), .CK(clock), .Q(
        decode_regfile_intregs_27__6_) );
  DFF_X2 decode_regfile_intregs_reg_27__7_ ( .D(n7083), .CK(clock), .Q(
        decode_regfile_intregs_27__7_) );
  DFF_X2 decode_regfile_intregs_reg_27__8_ ( .D(n7082), .CK(clock), .Q(
        decode_regfile_intregs_27__8_) );
  DFF_X2 decode_regfile_intregs_reg_27__9_ ( .D(n7081), .CK(clock), .Q(
        decode_regfile_intregs_27__9_) );
  DFF_X2 decode_regfile_intregs_reg_27__10_ ( .D(n7080), .CK(clock), .Q(
        decode_regfile_intregs_27__10_) );
  DFF_X2 decode_regfile_intregs_reg_27__11_ ( .D(n7079), .CK(clock), .Q(
        decode_regfile_intregs_27__11_) );
  DFF_X2 decode_regfile_intregs_reg_27__12_ ( .D(n7078), .CK(clock), .Q(
        decode_regfile_intregs_27__12_) );
  DFF_X2 decode_regfile_intregs_reg_27__13_ ( .D(n7077), .CK(clock), .Q(
        decode_regfile_intregs_27__13_) );
  DFF_X2 decode_regfile_intregs_reg_27__14_ ( .D(n7076), .CK(clock), .Q(
        decode_regfile_intregs_27__14_) );
  DFF_X2 decode_regfile_intregs_reg_27__15_ ( .D(n7075), .CK(clock), .Q(
        decode_regfile_intregs_27__15_) );
  DFF_X2 decode_regfile_intregs_reg_27__16_ ( .D(n7074), .CK(clock), .Q(
        decode_regfile_intregs_27__16_) );
  DFF_X2 decode_regfile_intregs_reg_27__17_ ( .D(n7073), .CK(clock), .Q(
        decode_regfile_intregs_27__17_) );
  DFF_X2 decode_regfile_intregs_reg_27__18_ ( .D(n7072), .CK(clock), .Q(
        decode_regfile_intregs_27__18_) );
  DFF_X2 decode_regfile_intregs_reg_27__19_ ( .D(n7071), .CK(clock), .Q(
        decode_regfile_intregs_27__19_) );
  DFF_X2 decode_regfile_intregs_reg_27__20_ ( .D(n7070), .CK(clock), .Q(
        decode_regfile_intregs_27__20_) );
  DFF_X2 decode_regfile_intregs_reg_27__21_ ( .D(n7069), .CK(clock), .Q(
        decode_regfile_intregs_27__21_) );
  DFF_X2 decode_regfile_intregs_reg_27__22_ ( .D(n7068), .CK(clock), .Q(
        decode_regfile_intregs_27__22_) );
  DFF_X2 decode_regfile_intregs_reg_27__23_ ( .D(n7067), .CK(clock), .Q(
        decode_regfile_intregs_27__23_) );
  DFF_X2 decode_regfile_intregs_reg_27__24_ ( .D(n7066), .CK(clock), .Q(
        decode_regfile_intregs_27__24_) );
  DFF_X2 decode_regfile_intregs_reg_27__25_ ( .D(n7065), .CK(clock), .Q(
        decode_regfile_intregs_27__25_) );
  DFF_X2 decode_regfile_intregs_reg_27__26_ ( .D(n7064), .CK(clock), .Q(
        decode_regfile_intregs_27__26_) );
  DFF_X2 decode_regfile_intregs_reg_27__27_ ( .D(n7063), .CK(clock), .Q(
        decode_regfile_intregs_27__27_) );
  DFF_X2 decode_regfile_intregs_reg_27__28_ ( .D(n7062), .CK(clock), .Q(
        decode_regfile_intregs_27__28_) );
  DFF_X2 decode_regfile_intregs_reg_27__29_ ( .D(n7061), .CK(clock), .Q(
        decode_regfile_intregs_27__29_) );
  DFF_X2 decode_regfile_intregs_reg_27__30_ ( .D(n7060), .CK(clock), .Q(
        decode_regfile_intregs_27__30_) );
  DFF_X2 decode_regfile_intregs_reg_27__31_ ( .D(n7059), .CK(clock), .Q(
        decode_regfile_intregs_27__31_) );
  DFF_X2 decode_regfile_intregs_reg_26__0_ ( .D(n7058), .CK(clock), .Q(
        decode_regfile_intregs_26__0_) );
  DFF_X2 decode_regfile_intregs_reg_26__1_ ( .D(n7057), .CK(clock), .Q(
        decode_regfile_intregs_26__1_) );
  DFF_X2 decode_regfile_intregs_reg_26__2_ ( .D(n7056), .CK(clock), .Q(
        decode_regfile_intregs_26__2_) );
  DFF_X2 decode_regfile_intregs_reg_26__3_ ( .D(n7055), .CK(clock), .Q(
        decode_regfile_intregs_26__3_) );
  DFF_X2 decode_regfile_intregs_reg_26__4_ ( .D(n7054), .CK(clock), .Q(
        decode_regfile_intregs_26__4_) );
  DFF_X2 decode_regfile_intregs_reg_26__5_ ( .D(n7053), .CK(clock), .Q(
        decode_regfile_intregs_26__5_) );
  DFF_X2 decode_regfile_intregs_reg_26__6_ ( .D(n7052), .CK(clock), .Q(
        decode_regfile_intregs_26__6_) );
  DFF_X2 decode_regfile_intregs_reg_26__7_ ( .D(n7051), .CK(clock), .Q(
        decode_regfile_intregs_26__7_) );
  DFF_X2 decode_regfile_intregs_reg_26__8_ ( .D(n7050), .CK(clock), .Q(
        decode_regfile_intregs_26__8_) );
  DFF_X2 decode_regfile_intregs_reg_26__9_ ( .D(n7049), .CK(clock), .Q(
        decode_regfile_intregs_26__9_) );
  DFF_X2 decode_regfile_intregs_reg_26__10_ ( .D(n7048), .CK(clock), .Q(
        decode_regfile_intregs_26__10_) );
  DFF_X2 decode_regfile_intregs_reg_26__11_ ( .D(n7047), .CK(clock), .Q(
        decode_regfile_intregs_26__11_) );
  DFF_X2 decode_regfile_intregs_reg_26__12_ ( .D(n7046), .CK(clock), .Q(
        decode_regfile_intregs_26__12_) );
  DFF_X2 decode_regfile_intregs_reg_26__13_ ( .D(n7045), .CK(clock), .Q(
        decode_regfile_intregs_26__13_) );
  DFF_X2 decode_regfile_intregs_reg_26__14_ ( .D(n7044), .CK(clock), .Q(
        decode_regfile_intregs_26__14_) );
  DFF_X2 decode_regfile_intregs_reg_26__15_ ( .D(n7043), .CK(clock), .Q(
        decode_regfile_intregs_26__15_) );
  DFF_X2 decode_regfile_intregs_reg_26__16_ ( .D(n7042), .CK(clock), .Q(
        decode_regfile_intregs_26__16_) );
  DFF_X2 decode_regfile_intregs_reg_26__17_ ( .D(n7041), .CK(clock), .Q(
        decode_regfile_intregs_26__17_) );
  DFF_X2 decode_regfile_intregs_reg_26__18_ ( .D(n7040), .CK(clock), .Q(
        decode_regfile_intregs_26__18_) );
  DFF_X2 decode_regfile_intregs_reg_26__19_ ( .D(n7039), .CK(clock), .Q(
        decode_regfile_intregs_26__19_) );
  DFF_X2 decode_regfile_intregs_reg_26__20_ ( .D(n7038), .CK(clock), .Q(
        decode_regfile_intregs_26__20_) );
  DFF_X2 decode_regfile_intregs_reg_26__21_ ( .D(n7037), .CK(clock), .Q(
        decode_regfile_intregs_26__21_) );
  DFF_X2 decode_regfile_intregs_reg_26__22_ ( .D(n7036), .CK(clock), .Q(
        decode_regfile_intregs_26__22_) );
  DFF_X2 decode_regfile_intregs_reg_26__23_ ( .D(n7035), .CK(clock), .Q(
        decode_regfile_intregs_26__23_) );
  DFF_X2 decode_regfile_intregs_reg_26__24_ ( .D(n7034), .CK(clock), .Q(
        decode_regfile_intregs_26__24_) );
  DFF_X2 decode_regfile_intregs_reg_26__25_ ( .D(n7033), .CK(clock), .Q(
        decode_regfile_intregs_26__25_) );
  DFF_X2 decode_regfile_intregs_reg_26__26_ ( .D(n7032), .CK(clock), .Q(
        decode_regfile_intregs_26__26_) );
  DFF_X2 decode_regfile_intregs_reg_26__27_ ( .D(n7031), .CK(clock), .Q(
        decode_regfile_intregs_26__27_) );
  DFF_X2 decode_regfile_intregs_reg_26__28_ ( .D(n7030), .CK(clock), .Q(
        decode_regfile_intregs_26__28_) );
  DFF_X2 decode_regfile_intregs_reg_26__29_ ( .D(n7029), .CK(clock), .Q(
        decode_regfile_intregs_26__29_) );
  DFF_X2 decode_regfile_intregs_reg_26__30_ ( .D(n7028), .CK(clock), .Q(
        decode_regfile_intregs_26__30_) );
  DFF_X2 decode_regfile_intregs_reg_26__31_ ( .D(n7027), .CK(clock), .Q(
        decode_regfile_intregs_26__31_) );
  DFF_X2 decode_regfile_intregs_reg_25__0_ ( .D(n7026), .CK(clock), .Q(
        decode_regfile_intregs_25__0_) );
  DFF_X2 decode_regfile_intregs_reg_25__1_ ( .D(n7025), .CK(clock), .Q(
        decode_regfile_intregs_25__1_) );
  DFF_X2 decode_regfile_intregs_reg_25__2_ ( .D(n7024), .CK(clock), .Q(
        decode_regfile_intregs_25__2_) );
  DFF_X2 decode_regfile_intregs_reg_25__3_ ( .D(n7023), .CK(clock), .Q(
        decode_regfile_intregs_25__3_) );
  DFF_X2 decode_regfile_intregs_reg_25__4_ ( .D(n7022), .CK(clock), .Q(
        decode_regfile_intregs_25__4_) );
  DFF_X2 decode_regfile_intregs_reg_25__5_ ( .D(n7021), .CK(clock), .Q(
        decode_regfile_intregs_25__5_) );
  DFF_X2 decode_regfile_intregs_reg_25__6_ ( .D(n7020), .CK(clock), .Q(
        decode_regfile_intregs_25__6_) );
  DFF_X2 decode_regfile_intregs_reg_25__7_ ( .D(n7019), .CK(clock), .Q(
        decode_regfile_intregs_25__7_) );
  DFF_X2 decode_regfile_intregs_reg_25__8_ ( .D(n7018), .CK(clock), .Q(
        decode_regfile_intregs_25__8_) );
  DFF_X2 decode_regfile_intregs_reg_25__9_ ( .D(n7017), .CK(clock), .Q(
        decode_regfile_intregs_25__9_) );
  DFF_X2 decode_regfile_intregs_reg_25__10_ ( .D(n7016), .CK(clock), .Q(
        decode_regfile_intregs_25__10_) );
  DFF_X2 decode_regfile_intregs_reg_25__11_ ( .D(n7015), .CK(clock), .Q(
        decode_regfile_intregs_25__11_) );
  DFF_X2 decode_regfile_intregs_reg_25__12_ ( .D(n7014), .CK(clock), .Q(
        decode_regfile_intregs_25__12_) );
  DFF_X2 decode_regfile_intregs_reg_25__13_ ( .D(n7013), .CK(clock), .Q(
        decode_regfile_intregs_25__13_) );
  DFF_X2 decode_regfile_intregs_reg_25__14_ ( .D(n7012), .CK(clock), .Q(
        decode_regfile_intregs_25__14_) );
  DFF_X2 decode_regfile_intregs_reg_25__15_ ( .D(n7011), .CK(clock), .Q(
        decode_regfile_intregs_25__15_) );
  DFF_X2 decode_regfile_intregs_reg_25__16_ ( .D(n7010), .CK(clock), .Q(
        decode_regfile_intregs_25__16_) );
  DFF_X2 decode_regfile_intregs_reg_25__17_ ( .D(n7009), .CK(clock), .Q(
        decode_regfile_intregs_25__17_) );
  DFF_X2 decode_regfile_intregs_reg_25__18_ ( .D(n7008), .CK(clock), .Q(
        decode_regfile_intregs_25__18_) );
  DFF_X2 decode_regfile_intregs_reg_25__19_ ( .D(n7007), .CK(clock), .Q(
        decode_regfile_intregs_25__19_) );
  DFF_X2 decode_regfile_intregs_reg_25__20_ ( .D(n7006), .CK(clock), .Q(
        decode_regfile_intregs_25__20_) );
  DFF_X2 decode_regfile_intregs_reg_25__21_ ( .D(n7005), .CK(clock), .Q(
        decode_regfile_intregs_25__21_) );
  DFF_X2 decode_regfile_intregs_reg_25__22_ ( .D(n7004), .CK(clock), .Q(
        decode_regfile_intregs_25__22_) );
  DFF_X2 decode_regfile_intregs_reg_25__23_ ( .D(n7003), .CK(clock), .Q(
        decode_regfile_intregs_25__23_) );
  DFF_X2 decode_regfile_intregs_reg_25__24_ ( .D(n7002), .CK(clock), .Q(
        decode_regfile_intregs_25__24_) );
  DFF_X2 decode_regfile_intregs_reg_25__25_ ( .D(n7001), .CK(clock), .Q(
        decode_regfile_intregs_25__25_) );
  DFF_X2 decode_regfile_intregs_reg_25__26_ ( .D(n7000), .CK(clock), .Q(
        decode_regfile_intregs_25__26_) );
  DFF_X2 decode_regfile_intregs_reg_25__27_ ( .D(n6999), .CK(clock), .Q(
        decode_regfile_intregs_25__27_) );
  DFF_X2 decode_regfile_intregs_reg_25__28_ ( .D(n6998), .CK(clock), .Q(
        decode_regfile_intregs_25__28_) );
  DFF_X2 decode_regfile_intregs_reg_25__29_ ( .D(n6997), .CK(clock), .Q(
        decode_regfile_intregs_25__29_) );
  DFF_X2 decode_regfile_intregs_reg_25__30_ ( .D(n6996), .CK(clock), .Q(
        decode_regfile_intregs_25__30_) );
  DFF_X2 decode_regfile_intregs_reg_25__31_ ( .D(n6995), .CK(clock), .Q(
        decode_regfile_intregs_25__31_) );
  DFF_X2 decode_regfile_intregs_reg_24__0_ ( .D(n6994), .CK(clock), .Q(
        decode_regfile_intregs_24__0_) );
  DFF_X2 decode_regfile_intregs_reg_24__1_ ( .D(n6993), .CK(clock), .Q(
        decode_regfile_intregs_24__1_) );
  DFF_X2 decode_regfile_intregs_reg_24__2_ ( .D(n6992), .CK(clock), .Q(
        decode_regfile_intregs_24__2_) );
  DFF_X2 decode_regfile_intregs_reg_24__3_ ( .D(n6991), .CK(clock), .Q(
        decode_regfile_intregs_24__3_) );
  DFF_X2 decode_regfile_intregs_reg_24__4_ ( .D(n6990), .CK(clock), .Q(
        decode_regfile_intregs_24__4_) );
  DFF_X2 decode_regfile_intregs_reg_24__5_ ( .D(n6989), .CK(clock), .Q(
        decode_regfile_intregs_24__5_) );
  DFF_X2 decode_regfile_intregs_reg_24__6_ ( .D(n6988), .CK(clock), .Q(
        decode_regfile_intregs_24__6_) );
  DFF_X2 decode_regfile_intregs_reg_24__7_ ( .D(n6987), .CK(clock), .Q(
        decode_regfile_intregs_24__7_) );
  DFF_X2 decode_regfile_intregs_reg_24__8_ ( .D(n6986), .CK(clock), .Q(
        decode_regfile_intregs_24__8_) );
  DFF_X2 decode_regfile_intregs_reg_24__9_ ( .D(n6985), .CK(clock), .Q(
        decode_regfile_intregs_24__9_) );
  DFF_X2 decode_regfile_intregs_reg_24__10_ ( .D(n6984), .CK(clock), .Q(
        decode_regfile_intregs_24__10_) );
  DFF_X2 decode_regfile_intregs_reg_24__11_ ( .D(n6983), .CK(clock), .Q(
        decode_regfile_intregs_24__11_) );
  DFF_X2 decode_regfile_intregs_reg_24__12_ ( .D(n6982), .CK(clock), .Q(
        decode_regfile_intregs_24__12_) );
  DFF_X2 decode_regfile_intregs_reg_24__13_ ( .D(n6981), .CK(clock), .Q(
        decode_regfile_intregs_24__13_) );
  DFF_X2 decode_regfile_intregs_reg_24__14_ ( .D(n6980), .CK(clock), .Q(
        decode_regfile_intregs_24__14_) );
  DFF_X2 decode_regfile_intregs_reg_24__15_ ( .D(n6979), .CK(clock), .Q(
        decode_regfile_intregs_24__15_) );
  DFF_X2 decode_regfile_intregs_reg_24__16_ ( .D(n6978), .CK(clock), .Q(
        decode_regfile_intregs_24__16_) );
  DFF_X2 decode_regfile_intregs_reg_24__17_ ( .D(n6977), .CK(clock), .Q(
        decode_regfile_intregs_24__17_) );
  DFF_X2 decode_regfile_intregs_reg_24__18_ ( .D(n6976), .CK(clock), .Q(
        decode_regfile_intregs_24__18_) );
  DFF_X2 decode_regfile_intregs_reg_24__19_ ( .D(n6975), .CK(clock), .Q(
        decode_regfile_intregs_24__19_) );
  DFF_X2 decode_regfile_intregs_reg_24__20_ ( .D(n6974), .CK(clock), .Q(
        decode_regfile_intregs_24__20_) );
  DFF_X2 decode_regfile_intregs_reg_24__21_ ( .D(n6973), .CK(clock), .Q(
        decode_regfile_intregs_24__21_) );
  DFF_X2 decode_regfile_intregs_reg_24__22_ ( .D(n6972), .CK(clock), .Q(
        decode_regfile_intregs_24__22_) );
  DFF_X2 decode_regfile_intregs_reg_24__23_ ( .D(n6971), .CK(clock), .Q(
        decode_regfile_intregs_24__23_) );
  DFF_X2 decode_regfile_intregs_reg_24__24_ ( .D(n6970), .CK(clock), .Q(
        decode_regfile_intregs_24__24_) );
  DFF_X2 decode_regfile_intregs_reg_24__25_ ( .D(n6969), .CK(clock), .Q(
        decode_regfile_intregs_24__25_) );
  DFF_X2 decode_regfile_intregs_reg_24__26_ ( .D(n6968), .CK(clock), .Q(
        decode_regfile_intregs_24__26_) );
  DFF_X2 decode_regfile_intregs_reg_24__27_ ( .D(n6967), .CK(clock), .Q(
        decode_regfile_intregs_24__27_) );
  DFF_X2 decode_regfile_intregs_reg_24__28_ ( .D(n6966), .CK(clock), .Q(
        decode_regfile_intregs_24__28_) );
  DFF_X2 decode_regfile_intregs_reg_24__29_ ( .D(n6965), .CK(clock), .Q(
        decode_regfile_intregs_24__29_) );
  DFF_X2 decode_regfile_intregs_reg_24__30_ ( .D(n6964), .CK(clock), .Q(
        decode_regfile_intregs_24__30_) );
  DFF_X2 decode_regfile_intregs_reg_24__31_ ( .D(n6963), .CK(clock), .Q(
        decode_regfile_intregs_24__31_) );
  DFF_X2 decode_regfile_intregs_reg_23__0_ ( .D(n6962), .CK(clock), .Q(
        decode_regfile_intregs_23__0_) );
  DFF_X2 decode_regfile_intregs_reg_23__1_ ( .D(n6961), .CK(clock), .Q(
        decode_regfile_intregs_23__1_) );
  DFF_X2 decode_regfile_intregs_reg_23__2_ ( .D(n6960), .CK(clock), .Q(
        decode_regfile_intregs_23__2_) );
  DFF_X2 decode_regfile_intregs_reg_23__3_ ( .D(n6959), .CK(clock), .Q(
        decode_regfile_intregs_23__3_) );
  DFF_X2 decode_regfile_intregs_reg_23__4_ ( .D(n6958), .CK(clock), .Q(
        decode_regfile_intregs_23__4_) );
  DFF_X2 decode_regfile_intregs_reg_23__5_ ( .D(n6957), .CK(clock), .Q(
        decode_regfile_intregs_23__5_) );
  DFF_X2 decode_regfile_intregs_reg_23__6_ ( .D(n6956), .CK(clock), .Q(
        decode_regfile_intregs_23__6_) );
  DFF_X2 decode_regfile_intregs_reg_23__7_ ( .D(n6955), .CK(clock), .Q(
        decode_regfile_intregs_23__7_) );
  DFF_X2 decode_regfile_intregs_reg_23__8_ ( .D(n6954), .CK(clock), .Q(
        decode_regfile_intregs_23__8_) );
  DFF_X2 decode_regfile_intregs_reg_23__9_ ( .D(n6953), .CK(clock), .Q(
        decode_regfile_intregs_23__9_) );
  DFF_X2 decode_regfile_intregs_reg_23__10_ ( .D(n6952), .CK(clock), .Q(
        decode_regfile_intregs_23__10_) );
  DFF_X2 decode_regfile_intregs_reg_23__11_ ( .D(n6951), .CK(clock), .Q(
        decode_regfile_intregs_23__11_) );
  DFF_X2 decode_regfile_intregs_reg_23__12_ ( .D(n6950), .CK(clock), .Q(
        decode_regfile_intregs_23__12_) );
  DFF_X2 decode_regfile_intregs_reg_23__13_ ( .D(n6949), .CK(clock), .Q(
        decode_regfile_intregs_23__13_) );
  DFF_X2 decode_regfile_intregs_reg_23__14_ ( .D(n6948), .CK(clock), .Q(
        decode_regfile_intregs_23__14_) );
  DFF_X2 decode_regfile_intregs_reg_23__15_ ( .D(n6947), .CK(clock), .Q(
        decode_regfile_intregs_23__15_) );
  DFF_X2 decode_regfile_intregs_reg_23__16_ ( .D(n6946), .CK(clock), .Q(
        decode_regfile_intregs_23__16_) );
  DFF_X2 decode_regfile_intregs_reg_23__17_ ( .D(n6945), .CK(clock), .Q(
        decode_regfile_intregs_23__17_) );
  DFF_X2 decode_regfile_intregs_reg_23__18_ ( .D(n6944), .CK(clock), .Q(
        decode_regfile_intregs_23__18_) );
  DFF_X2 decode_regfile_intregs_reg_23__19_ ( .D(n6943), .CK(clock), .Q(
        decode_regfile_intregs_23__19_) );
  DFF_X2 decode_regfile_intregs_reg_23__20_ ( .D(n6942), .CK(clock), .Q(
        decode_regfile_intregs_23__20_) );
  DFF_X2 decode_regfile_intregs_reg_23__21_ ( .D(n6941), .CK(clock), .Q(
        decode_regfile_intregs_23__21_) );
  DFF_X2 decode_regfile_intregs_reg_23__22_ ( .D(n6940), .CK(clock), .Q(
        decode_regfile_intregs_23__22_) );
  DFF_X2 decode_regfile_intregs_reg_23__23_ ( .D(n6939), .CK(clock), .Q(
        decode_regfile_intregs_23__23_) );
  DFF_X2 decode_regfile_intregs_reg_23__24_ ( .D(n6938), .CK(clock), .Q(
        decode_regfile_intregs_23__24_) );
  DFF_X2 decode_regfile_intregs_reg_23__25_ ( .D(n6937), .CK(clock), .Q(
        decode_regfile_intregs_23__25_) );
  DFF_X2 decode_regfile_intregs_reg_23__26_ ( .D(n6936), .CK(clock), .Q(
        decode_regfile_intregs_23__26_) );
  DFF_X2 decode_regfile_intregs_reg_23__27_ ( .D(n6935), .CK(clock), .Q(
        decode_regfile_intregs_23__27_) );
  DFF_X2 decode_regfile_intregs_reg_23__28_ ( .D(n6934), .CK(clock), .Q(
        decode_regfile_intregs_23__28_) );
  DFF_X2 decode_regfile_intregs_reg_23__29_ ( .D(n6933), .CK(clock), .Q(
        decode_regfile_intregs_23__29_) );
  DFF_X2 decode_regfile_intregs_reg_23__30_ ( .D(n6932), .CK(clock), .Q(
        decode_regfile_intregs_23__30_) );
  DFF_X2 decode_regfile_intregs_reg_23__31_ ( .D(n6931), .CK(clock), .Q(
        decode_regfile_intregs_23__31_) );
  DFF_X2 decode_regfile_intregs_reg_22__0_ ( .D(n6930), .CK(clock), .Q(
        decode_regfile_intregs_22__0_) );
  DFF_X2 decode_regfile_intregs_reg_22__1_ ( .D(n6929), .CK(clock), .Q(
        decode_regfile_intregs_22__1_) );
  DFF_X2 decode_regfile_intregs_reg_22__2_ ( .D(n6928), .CK(clock), .Q(
        decode_regfile_intregs_22__2_) );
  DFF_X2 decode_regfile_intregs_reg_22__3_ ( .D(n6927), .CK(clock), .Q(
        decode_regfile_intregs_22__3_) );
  DFF_X2 decode_regfile_intregs_reg_22__4_ ( .D(n6926), .CK(clock), .Q(
        decode_regfile_intregs_22__4_) );
  DFF_X2 decode_regfile_intregs_reg_22__5_ ( .D(n6925), .CK(clock), .Q(
        decode_regfile_intregs_22__5_) );
  DFF_X2 decode_regfile_intregs_reg_22__6_ ( .D(n6924), .CK(clock), .Q(
        decode_regfile_intregs_22__6_) );
  DFF_X2 decode_regfile_intregs_reg_22__7_ ( .D(n6923), .CK(clock), .Q(
        decode_regfile_intregs_22__7_) );
  DFF_X2 decode_regfile_intregs_reg_22__8_ ( .D(n6922), .CK(clock), .Q(
        decode_regfile_intregs_22__8_) );
  DFF_X2 decode_regfile_intregs_reg_22__9_ ( .D(n6921), .CK(clock), .Q(
        decode_regfile_intregs_22__9_) );
  DFF_X2 decode_regfile_intregs_reg_22__10_ ( .D(n6920), .CK(clock), .Q(
        decode_regfile_intregs_22__10_) );
  DFF_X2 decode_regfile_intregs_reg_22__11_ ( .D(n6919), .CK(clock), .Q(
        decode_regfile_intregs_22__11_) );
  DFF_X2 decode_regfile_intregs_reg_22__12_ ( .D(n6918), .CK(clock), .Q(
        decode_regfile_intregs_22__12_) );
  DFF_X2 decode_regfile_intregs_reg_22__13_ ( .D(n6917), .CK(clock), .Q(
        decode_regfile_intregs_22__13_) );
  DFF_X2 decode_regfile_intregs_reg_22__14_ ( .D(n6916), .CK(clock), .Q(
        decode_regfile_intregs_22__14_) );
  DFF_X2 decode_regfile_intregs_reg_22__15_ ( .D(n6915), .CK(clock), .Q(
        decode_regfile_intregs_22__15_) );
  DFF_X2 decode_regfile_intregs_reg_22__16_ ( .D(n6914), .CK(clock), .Q(
        decode_regfile_intregs_22__16_) );
  DFF_X2 decode_regfile_intregs_reg_22__17_ ( .D(n6913), .CK(clock), .Q(
        decode_regfile_intregs_22__17_) );
  DFF_X2 decode_regfile_intregs_reg_22__18_ ( .D(n6912), .CK(clock), .Q(
        decode_regfile_intregs_22__18_) );
  DFF_X2 decode_regfile_intregs_reg_22__19_ ( .D(n6911), .CK(clock), .Q(
        decode_regfile_intregs_22__19_) );
  DFF_X2 decode_regfile_intregs_reg_22__20_ ( .D(n6910), .CK(clock), .Q(
        decode_regfile_intregs_22__20_) );
  DFF_X2 decode_regfile_intregs_reg_22__21_ ( .D(n6909), .CK(clock), .Q(
        decode_regfile_intregs_22__21_) );
  DFF_X2 decode_regfile_intregs_reg_22__22_ ( .D(n6908), .CK(clock), .Q(
        decode_regfile_intregs_22__22_) );
  DFF_X2 decode_regfile_intregs_reg_22__23_ ( .D(n6907), .CK(clock), .Q(
        decode_regfile_intregs_22__23_) );
  DFF_X2 decode_regfile_intregs_reg_22__24_ ( .D(n6906), .CK(clock), .Q(
        decode_regfile_intregs_22__24_) );
  DFF_X2 decode_regfile_intregs_reg_22__25_ ( .D(n6905), .CK(clock), .Q(
        decode_regfile_intregs_22__25_) );
  DFF_X2 decode_regfile_intregs_reg_22__26_ ( .D(n6904), .CK(clock), .Q(
        decode_regfile_intregs_22__26_) );
  DFF_X2 decode_regfile_intregs_reg_22__27_ ( .D(n6903), .CK(clock), .Q(
        decode_regfile_intregs_22__27_) );
  DFF_X2 decode_regfile_intregs_reg_22__28_ ( .D(n6902), .CK(clock), .Q(
        decode_regfile_intregs_22__28_) );
  DFF_X2 decode_regfile_intregs_reg_22__29_ ( .D(n6901), .CK(clock), .Q(
        decode_regfile_intregs_22__29_) );
  DFF_X2 decode_regfile_intregs_reg_22__30_ ( .D(n6900), .CK(clock), .Q(
        decode_regfile_intregs_22__30_) );
  DFF_X2 decode_regfile_intregs_reg_22__31_ ( .D(n6899), .CK(clock), .Q(
        decode_regfile_intregs_22__31_) );
  DFF_X2 decode_regfile_intregs_reg_21__0_ ( .D(n6898), .CK(clock), .Q(
        decode_regfile_intregs_21__0_) );
  DFF_X2 decode_regfile_intregs_reg_21__1_ ( .D(n6897), .CK(clock), .Q(
        decode_regfile_intregs_21__1_) );
  DFF_X2 decode_regfile_intregs_reg_21__2_ ( .D(n6896), .CK(clock), .Q(
        decode_regfile_intregs_21__2_) );
  DFF_X2 decode_regfile_intregs_reg_21__3_ ( .D(n6895), .CK(clock), .Q(
        decode_regfile_intregs_21__3_) );
  DFF_X2 decode_regfile_intregs_reg_21__4_ ( .D(n6894), .CK(clock), .Q(
        decode_regfile_intregs_21__4_) );
  DFF_X2 decode_regfile_intregs_reg_21__5_ ( .D(n6893), .CK(clock), .Q(
        decode_regfile_intregs_21__5_) );
  DFF_X2 decode_regfile_intregs_reg_21__6_ ( .D(n6892), .CK(clock), .Q(
        decode_regfile_intregs_21__6_) );
  DFF_X2 decode_regfile_intregs_reg_21__7_ ( .D(n6891), .CK(clock), .Q(
        decode_regfile_intregs_21__7_) );
  DFF_X2 decode_regfile_intregs_reg_21__8_ ( .D(n6890), .CK(clock), .Q(
        decode_regfile_intregs_21__8_) );
  DFF_X2 decode_regfile_intregs_reg_21__9_ ( .D(n6889), .CK(clock), .Q(
        decode_regfile_intregs_21__9_) );
  DFF_X2 decode_regfile_intregs_reg_21__10_ ( .D(n6888), .CK(clock), .Q(
        decode_regfile_intregs_21__10_) );
  DFF_X2 decode_regfile_intregs_reg_21__11_ ( .D(n6887), .CK(clock), .Q(
        decode_regfile_intregs_21__11_) );
  DFF_X2 decode_regfile_intregs_reg_21__12_ ( .D(n6886), .CK(clock), .Q(
        decode_regfile_intregs_21__12_) );
  DFF_X2 decode_regfile_intregs_reg_21__13_ ( .D(n6885), .CK(clock), .Q(
        decode_regfile_intregs_21__13_) );
  DFF_X2 decode_regfile_intregs_reg_21__14_ ( .D(n6884), .CK(clock), .Q(
        decode_regfile_intregs_21__14_) );
  DFF_X2 decode_regfile_intregs_reg_21__15_ ( .D(n6883), .CK(clock), .Q(
        decode_regfile_intregs_21__15_) );
  DFF_X2 decode_regfile_intregs_reg_21__16_ ( .D(n6882), .CK(clock), .Q(
        decode_regfile_intregs_21__16_) );
  DFF_X2 decode_regfile_intregs_reg_21__17_ ( .D(n6881), .CK(clock), .Q(
        decode_regfile_intregs_21__17_) );
  DFF_X2 decode_regfile_intregs_reg_21__18_ ( .D(n6880), .CK(clock), .Q(
        decode_regfile_intregs_21__18_) );
  DFF_X2 decode_regfile_intregs_reg_21__19_ ( .D(n6879), .CK(clock), .Q(
        decode_regfile_intregs_21__19_) );
  DFF_X2 decode_regfile_intregs_reg_21__20_ ( .D(n6878), .CK(clock), .Q(
        decode_regfile_intregs_21__20_) );
  DFF_X2 decode_regfile_intregs_reg_21__21_ ( .D(n6877), .CK(clock), .Q(
        decode_regfile_intregs_21__21_) );
  DFF_X2 decode_regfile_intregs_reg_21__22_ ( .D(n6876), .CK(clock), .Q(
        decode_regfile_intregs_21__22_) );
  DFF_X2 decode_regfile_intregs_reg_21__23_ ( .D(n6875), .CK(clock), .Q(
        decode_regfile_intregs_21__23_) );
  DFF_X2 decode_regfile_intregs_reg_21__24_ ( .D(n6874), .CK(clock), .Q(
        decode_regfile_intregs_21__24_) );
  DFF_X2 decode_regfile_intregs_reg_21__25_ ( .D(n6873), .CK(clock), .Q(
        decode_regfile_intregs_21__25_) );
  DFF_X2 decode_regfile_intregs_reg_21__26_ ( .D(n6872), .CK(clock), .Q(
        decode_regfile_intregs_21__26_) );
  DFF_X2 decode_regfile_intregs_reg_21__27_ ( .D(n6871), .CK(clock), .Q(
        decode_regfile_intregs_21__27_) );
  DFF_X2 decode_regfile_intregs_reg_21__28_ ( .D(n6870), .CK(clock), .Q(
        decode_regfile_intregs_21__28_) );
  DFF_X2 decode_regfile_intregs_reg_21__29_ ( .D(n6869), .CK(clock), .Q(
        decode_regfile_intregs_21__29_) );
  DFF_X2 decode_regfile_intregs_reg_21__30_ ( .D(n6868), .CK(clock), .Q(
        decode_regfile_intregs_21__30_) );
  DFF_X2 decode_regfile_intregs_reg_21__31_ ( .D(n6867), .CK(clock), .Q(
        decode_regfile_intregs_21__31_) );
  DFF_X2 decode_regfile_intregs_reg_20__0_ ( .D(n6866), .CK(clock), .Q(
        decode_regfile_intregs_20__0_) );
  DFF_X2 decode_regfile_intregs_reg_20__1_ ( .D(n6865), .CK(clock), .Q(
        decode_regfile_intregs_20__1_) );
  DFF_X2 decode_regfile_intregs_reg_20__2_ ( .D(n6864), .CK(clock), .Q(
        decode_regfile_intregs_20__2_) );
  DFF_X2 decode_regfile_intregs_reg_20__3_ ( .D(n6863), .CK(clock), .Q(
        decode_regfile_intregs_20__3_) );
  DFF_X2 decode_regfile_intregs_reg_20__4_ ( .D(n6862), .CK(clock), .Q(
        decode_regfile_intregs_20__4_) );
  DFF_X2 decode_regfile_intregs_reg_20__5_ ( .D(n6861), .CK(clock), .Q(
        decode_regfile_intregs_20__5_) );
  DFF_X2 decode_regfile_intregs_reg_20__6_ ( .D(n6860), .CK(clock), .Q(
        decode_regfile_intregs_20__6_) );
  DFF_X2 decode_regfile_intregs_reg_20__7_ ( .D(n6859), .CK(clock), .Q(
        decode_regfile_intregs_20__7_) );
  DFF_X2 decode_regfile_intregs_reg_20__8_ ( .D(n6858), .CK(clock), .Q(
        decode_regfile_intregs_20__8_) );
  DFF_X2 decode_regfile_intregs_reg_20__9_ ( .D(n6857), .CK(clock), .Q(
        decode_regfile_intregs_20__9_) );
  DFF_X2 decode_regfile_intregs_reg_20__10_ ( .D(n6856), .CK(clock), .Q(
        decode_regfile_intregs_20__10_) );
  DFF_X2 decode_regfile_intregs_reg_20__11_ ( .D(n6855), .CK(clock), .Q(
        decode_regfile_intregs_20__11_) );
  DFF_X2 decode_regfile_intregs_reg_20__12_ ( .D(n6854), .CK(clock), .Q(
        decode_regfile_intregs_20__12_) );
  DFF_X2 decode_regfile_intregs_reg_20__13_ ( .D(n6853), .CK(clock), .Q(
        decode_regfile_intregs_20__13_) );
  DFF_X2 decode_regfile_intregs_reg_20__14_ ( .D(n6852), .CK(clock), .Q(
        decode_regfile_intregs_20__14_) );
  DFF_X2 decode_regfile_intregs_reg_20__15_ ( .D(n6851), .CK(clock), .Q(
        decode_regfile_intregs_20__15_) );
  DFF_X2 decode_regfile_intregs_reg_20__16_ ( .D(n6850), .CK(clock), .Q(
        decode_regfile_intregs_20__16_) );
  DFF_X2 decode_regfile_intregs_reg_20__17_ ( .D(n6849), .CK(clock), .Q(
        decode_regfile_intregs_20__17_) );
  DFF_X2 decode_regfile_intregs_reg_20__18_ ( .D(n6848), .CK(clock), .Q(
        decode_regfile_intregs_20__18_) );
  DFF_X2 decode_regfile_intregs_reg_20__19_ ( .D(n6847), .CK(clock), .Q(
        decode_regfile_intregs_20__19_) );
  DFF_X2 decode_regfile_intregs_reg_20__20_ ( .D(n6846), .CK(clock), .Q(
        decode_regfile_intregs_20__20_) );
  DFF_X2 decode_regfile_intregs_reg_20__21_ ( .D(n6845), .CK(clock), .Q(
        decode_regfile_intregs_20__21_) );
  DFF_X2 decode_regfile_intregs_reg_20__22_ ( .D(n6844), .CK(clock), .Q(
        decode_regfile_intregs_20__22_) );
  DFF_X2 decode_regfile_intregs_reg_20__23_ ( .D(n6843), .CK(clock), .Q(
        decode_regfile_intregs_20__23_) );
  DFF_X2 decode_regfile_intregs_reg_20__24_ ( .D(n6842), .CK(clock), .Q(
        decode_regfile_intregs_20__24_) );
  DFF_X2 decode_regfile_intregs_reg_20__25_ ( .D(n6841), .CK(clock), .Q(
        decode_regfile_intregs_20__25_) );
  DFF_X2 decode_regfile_intregs_reg_20__26_ ( .D(n6840), .CK(clock), .Q(
        decode_regfile_intregs_20__26_) );
  DFF_X2 decode_regfile_intregs_reg_20__27_ ( .D(n6839), .CK(clock), .Q(
        decode_regfile_intregs_20__27_) );
  DFF_X2 decode_regfile_intregs_reg_20__28_ ( .D(n6838), .CK(clock), .Q(
        decode_regfile_intregs_20__28_) );
  DFF_X2 decode_regfile_intregs_reg_20__29_ ( .D(n6837), .CK(clock), .Q(
        decode_regfile_intregs_20__29_) );
  DFF_X2 decode_regfile_intregs_reg_20__30_ ( .D(n6836), .CK(clock), .Q(
        decode_regfile_intregs_20__30_) );
  DFF_X2 decode_regfile_intregs_reg_20__31_ ( .D(n6835), .CK(clock), .Q(
        decode_regfile_intregs_20__31_) );
  DFF_X2 decode_regfile_intregs_reg_19__0_ ( .D(n6834), .CK(clock), .Q(
        decode_regfile_intregs_19__0_) );
  DFF_X2 decode_regfile_intregs_reg_19__1_ ( .D(n6833), .CK(clock), .Q(
        decode_regfile_intregs_19__1_) );
  DFF_X2 decode_regfile_intregs_reg_19__2_ ( .D(n6832), .CK(clock), .Q(
        decode_regfile_intregs_19__2_) );
  DFF_X2 decode_regfile_intregs_reg_19__3_ ( .D(n6831), .CK(clock), .Q(
        decode_regfile_intregs_19__3_) );
  DFF_X2 decode_regfile_intregs_reg_19__4_ ( .D(n6830), .CK(clock), .Q(
        decode_regfile_intregs_19__4_) );
  DFF_X2 decode_regfile_intregs_reg_19__5_ ( .D(n6829), .CK(clock), .Q(
        decode_regfile_intregs_19__5_) );
  DFF_X2 decode_regfile_intregs_reg_19__6_ ( .D(n6828), .CK(clock), .Q(
        decode_regfile_intregs_19__6_) );
  DFF_X2 decode_regfile_intregs_reg_19__7_ ( .D(n6827), .CK(clock), .Q(
        decode_regfile_intregs_19__7_) );
  DFF_X2 decode_regfile_intregs_reg_19__8_ ( .D(n6826), .CK(clock), .Q(
        decode_regfile_intregs_19__8_) );
  DFF_X2 decode_regfile_intregs_reg_19__9_ ( .D(n6825), .CK(clock), .Q(
        decode_regfile_intregs_19__9_) );
  DFF_X2 decode_regfile_intregs_reg_19__10_ ( .D(n6824), .CK(clock), .Q(
        decode_regfile_intregs_19__10_) );
  DFF_X2 decode_regfile_intregs_reg_19__11_ ( .D(n6823), .CK(clock), .Q(
        decode_regfile_intregs_19__11_) );
  DFF_X2 decode_regfile_intregs_reg_19__12_ ( .D(n6822), .CK(clock), .Q(
        decode_regfile_intregs_19__12_) );
  DFF_X2 decode_regfile_intregs_reg_19__13_ ( .D(n6821), .CK(clock), .Q(
        decode_regfile_intregs_19__13_) );
  DFF_X2 decode_regfile_intregs_reg_19__14_ ( .D(n6820), .CK(clock), .Q(
        decode_regfile_intregs_19__14_) );
  DFF_X2 decode_regfile_intregs_reg_19__15_ ( .D(n6819), .CK(clock), .Q(
        decode_regfile_intregs_19__15_) );
  DFF_X2 decode_regfile_intregs_reg_19__16_ ( .D(n6818), .CK(clock), .Q(
        decode_regfile_intregs_19__16_) );
  DFF_X2 decode_regfile_intregs_reg_19__17_ ( .D(n6817), .CK(clock), .Q(
        decode_regfile_intregs_19__17_) );
  DFF_X2 decode_regfile_intregs_reg_19__18_ ( .D(n6816), .CK(clock), .Q(
        decode_regfile_intregs_19__18_) );
  DFF_X2 decode_regfile_intregs_reg_19__19_ ( .D(n6815), .CK(clock), .Q(
        decode_regfile_intregs_19__19_) );
  DFF_X2 decode_regfile_intregs_reg_19__20_ ( .D(n6814), .CK(clock), .Q(
        decode_regfile_intregs_19__20_) );
  DFF_X2 decode_regfile_intregs_reg_19__21_ ( .D(n6813), .CK(clock), .Q(
        decode_regfile_intregs_19__21_) );
  DFF_X2 decode_regfile_intregs_reg_19__22_ ( .D(n6812), .CK(clock), .Q(
        decode_regfile_intregs_19__22_) );
  DFF_X2 decode_regfile_intregs_reg_19__23_ ( .D(n6811), .CK(clock), .Q(
        decode_regfile_intregs_19__23_) );
  DFF_X2 decode_regfile_intregs_reg_19__24_ ( .D(n6810), .CK(clock), .Q(
        decode_regfile_intregs_19__24_) );
  DFF_X2 decode_regfile_intregs_reg_19__25_ ( .D(n6809), .CK(clock), .Q(
        decode_regfile_intregs_19__25_) );
  DFF_X2 decode_regfile_intregs_reg_19__26_ ( .D(n6808), .CK(clock), .Q(
        decode_regfile_intregs_19__26_) );
  DFF_X2 decode_regfile_intregs_reg_19__27_ ( .D(n6807), .CK(clock), .Q(
        decode_regfile_intregs_19__27_) );
  DFF_X2 decode_regfile_intregs_reg_19__28_ ( .D(n6806), .CK(clock), .Q(
        decode_regfile_intregs_19__28_) );
  DFF_X2 decode_regfile_intregs_reg_19__29_ ( .D(n6805), .CK(clock), .Q(
        decode_regfile_intregs_19__29_) );
  DFF_X2 decode_regfile_intregs_reg_19__30_ ( .D(n6804), .CK(clock), .Q(
        decode_regfile_intregs_19__30_) );
  DFF_X2 decode_regfile_intregs_reg_19__31_ ( .D(n6803), .CK(clock), .Q(
        decode_regfile_intregs_19__31_) );
  DFF_X2 decode_regfile_intregs_reg_18__0_ ( .D(n6802), .CK(clock), .Q(
        decode_regfile_intregs_18__0_) );
  DFF_X2 decode_regfile_intregs_reg_18__1_ ( .D(n6801), .CK(clock), .Q(
        decode_regfile_intregs_18__1_) );
  DFF_X2 decode_regfile_intregs_reg_18__2_ ( .D(n6800), .CK(clock), .Q(
        decode_regfile_intregs_18__2_) );
  DFF_X2 decode_regfile_intregs_reg_18__3_ ( .D(n6799), .CK(clock), .Q(
        decode_regfile_intregs_18__3_) );
  DFF_X2 decode_regfile_intregs_reg_18__4_ ( .D(n6798), .CK(clock), .Q(
        decode_regfile_intregs_18__4_) );
  DFF_X2 decode_regfile_intregs_reg_18__5_ ( .D(n6797), .CK(clock), .Q(
        decode_regfile_intregs_18__5_) );
  DFF_X2 decode_regfile_intregs_reg_18__6_ ( .D(n6796), .CK(clock), .Q(
        decode_regfile_intregs_18__6_) );
  DFF_X2 decode_regfile_intregs_reg_18__7_ ( .D(n6795), .CK(clock), .Q(
        decode_regfile_intregs_18__7_) );
  DFF_X2 decode_regfile_intregs_reg_18__8_ ( .D(n6794), .CK(clock), .Q(
        decode_regfile_intregs_18__8_) );
  DFF_X2 decode_regfile_intregs_reg_18__9_ ( .D(n6793), .CK(clock), .Q(
        decode_regfile_intregs_18__9_) );
  DFF_X2 decode_regfile_intregs_reg_18__10_ ( .D(n6792), .CK(clock), .Q(
        decode_regfile_intregs_18__10_) );
  DFF_X2 decode_regfile_intregs_reg_18__11_ ( .D(n6791), .CK(clock), .Q(
        decode_regfile_intregs_18__11_) );
  DFF_X2 decode_regfile_intregs_reg_18__12_ ( .D(n6790), .CK(clock), .Q(
        decode_regfile_intregs_18__12_) );
  DFF_X2 decode_regfile_intregs_reg_18__13_ ( .D(n6789), .CK(clock), .Q(
        decode_regfile_intregs_18__13_) );
  DFF_X2 decode_regfile_intregs_reg_18__14_ ( .D(n6788), .CK(clock), .Q(
        decode_regfile_intregs_18__14_) );
  DFF_X2 decode_regfile_intregs_reg_18__15_ ( .D(n6787), .CK(clock), .Q(
        decode_regfile_intregs_18__15_) );
  DFF_X2 decode_regfile_intregs_reg_18__16_ ( .D(n6786), .CK(clock), .Q(
        decode_regfile_intregs_18__16_) );
  DFF_X2 decode_regfile_intregs_reg_18__17_ ( .D(n6785), .CK(clock), .Q(
        decode_regfile_intregs_18__17_) );
  DFF_X2 decode_regfile_intregs_reg_18__18_ ( .D(n6784), .CK(clock), .Q(
        decode_regfile_intregs_18__18_) );
  DFF_X2 decode_regfile_intregs_reg_18__19_ ( .D(n6783), .CK(clock), .Q(
        decode_regfile_intregs_18__19_) );
  DFF_X2 decode_regfile_intregs_reg_18__20_ ( .D(n6782), .CK(clock), .Q(
        decode_regfile_intregs_18__20_) );
  DFF_X2 decode_regfile_intregs_reg_18__21_ ( .D(n6781), .CK(clock), .Q(
        decode_regfile_intregs_18__21_) );
  DFF_X2 decode_regfile_intregs_reg_18__22_ ( .D(n6780), .CK(clock), .Q(
        decode_regfile_intregs_18__22_) );
  DFF_X2 decode_regfile_intregs_reg_18__23_ ( .D(n6779), .CK(clock), .Q(
        decode_regfile_intregs_18__23_) );
  DFF_X2 decode_regfile_intregs_reg_18__24_ ( .D(n6778), .CK(clock), .Q(
        decode_regfile_intregs_18__24_) );
  DFF_X2 decode_regfile_intregs_reg_18__25_ ( .D(n6777), .CK(clock), .Q(
        decode_regfile_intregs_18__25_) );
  DFF_X2 decode_regfile_intregs_reg_18__26_ ( .D(n6776), .CK(clock), .Q(
        decode_regfile_intregs_18__26_) );
  DFF_X2 decode_regfile_intregs_reg_18__27_ ( .D(n6775), .CK(clock), .Q(
        decode_regfile_intregs_18__27_) );
  DFF_X2 decode_regfile_intregs_reg_18__28_ ( .D(n6774), .CK(clock), .Q(
        decode_regfile_intregs_18__28_) );
  DFF_X2 decode_regfile_intregs_reg_18__29_ ( .D(n6773), .CK(clock), .Q(
        decode_regfile_intregs_18__29_) );
  DFF_X2 decode_regfile_intregs_reg_18__30_ ( .D(n6772), .CK(clock), .Q(
        decode_regfile_intregs_18__30_) );
  DFF_X2 decode_regfile_intregs_reg_18__31_ ( .D(n6771), .CK(clock), .Q(
        decode_regfile_intregs_18__31_) );
  DFF_X2 decode_regfile_intregs_reg_17__0_ ( .D(n6770), .CK(clock), .Q(
        decode_regfile_intregs_17__0_) );
  DFF_X2 decode_regfile_intregs_reg_17__1_ ( .D(n6769), .CK(clock), .Q(
        decode_regfile_intregs_17__1_) );
  DFF_X2 decode_regfile_intregs_reg_17__2_ ( .D(n6768), .CK(clock), .Q(
        decode_regfile_intregs_17__2_) );
  DFF_X2 decode_regfile_intregs_reg_17__3_ ( .D(n6767), .CK(clock), .Q(
        decode_regfile_intregs_17__3_) );
  DFF_X2 decode_regfile_intregs_reg_17__4_ ( .D(n6766), .CK(clock), .Q(
        decode_regfile_intregs_17__4_) );
  DFF_X2 decode_regfile_intregs_reg_17__5_ ( .D(n6765), .CK(clock), .Q(
        decode_regfile_intregs_17__5_) );
  DFF_X2 decode_regfile_intregs_reg_17__6_ ( .D(n6764), .CK(clock), .Q(
        decode_regfile_intregs_17__6_) );
  DFF_X2 decode_regfile_intregs_reg_17__7_ ( .D(n6763), .CK(clock), .Q(
        decode_regfile_intregs_17__7_) );
  DFF_X2 decode_regfile_intregs_reg_17__8_ ( .D(n6762), .CK(clock), .Q(
        decode_regfile_intregs_17__8_) );
  DFF_X2 decode_regfile_intregs_reg_17__9_ ( .D(n6761), .CK(clock), .Q(
        decode_regfile_intregs_17__9_) );
  DFF_X2 decode_regfile_intregs_reg_17__10_ ( .D(n6760), .CK(clock), .Q(
        decode_regfile_intregs_17__10_) );
  DFF_X2 decode_regfile_intregs_reg_17__11_ ( .D(n6759), .CK(clock), .Q(
        decode_regfile_intregs_17__11_) );
  DFF_X2 decode_regfile_intregs_reg_17__12_ ( .D(n6758), .CK(clock), .Q(
        decode_regfile_intregs_17__12_) );
  DFF_X2 decode_regfile_intregs_reg_17__13_ ( .D(n6757), .CK(clock), .Q(
        decode_regfile_intregs_17__13_) );
  DFF_X2 decode_regfile_intregs_reg_17__14_ ( .D(n6756), .CK(clock), .Q(
        decode_regfile_intregs_17__14_) );
  DFF_X2 decode_regfile_intregs_reg_17__15_ ( .D(n6755), .CK(clock), .Q(
        decode_regfile_intregs_17__15_) );
  DFF_X2 decode_regfile_intregs_reg_17__16_ ( .D(n6754), .CK(clock), .Q(
        decode_regfile_intregs_17__16_) );
  DFF_X2 decode_regfile_intregs_reg_17__17_ ( .D(n6753), .CK(clock), .Q(
        decode_regfile_intregs_17__17_) );
  DFF_X2 decode_regfile_intregs_reg_17__18_ ( .D(n6752), .CK(clock), .Q(
        decode_regfile_intregs_17__18_) );
  DFF_X2 decode_regfile_intregs_reg_17__19_ ( .D(n6751), .CK(clock), .Q(
        decode_regfile_intregs_17__19_) );
  DFF_X2 decode_regfile_intregs_reg_17__20_ ( .D(n6750), .CK(clock), .Q(
        decode_regfile_intregs_17__20_) );
  DFF_X2 decode_regfile_intregs_reg_17__21_ ( .D(n6749), .CK(clock), .Q(
        decode_regfile_intregs_17__21_) );
  DFF_X2 decode_regfile_intregs_reg_17__22_ ( .D(n6748), .CK(clock), .Q(
        decode_regfile_intregs_17__22_) );
  DFF_X2 decode_regfile_intregs_reg_17__23_ ( .D(n6747), .CK(clock), .Q(
        decode_regfile_intregs_17__23_) );
  DFF_X2 decode_regfile_intregs_reg_17__24_ ( .D(n6746), .CK(clock), .Q(
        decode_regfile_intregs_17__24_) );
  DFF_X2 decode_regfile_intregs_reg_17__25_ ( .D(n6745), .CK(clock), .Q(
        decode_regfile_intregs_17__25_) );
  DFF_X2 decode_regfile_intregs_reg_17__26_ ( .D(n6744), .CK(clock), .Q(
        decode_regfile_intregs_17__26_) );
  DFF_X2 decode_regfile_intregs_reg_17__27_ ( .D(n6743), .CK(clock), .Q(
        decode_regfile_intregs_17__27_) );
  DFF_X2 decode_regfile_intregs_reg_17__28_ ( .D(n6742), .CK(clock), .Q(
        decode_regfile_intregs_17__28_) );
  DFF_X2 decode_regfile_intregs_reg_17__29_ ( .D(n6741), .CK(clock), .Q(
        decode_regfile_intregs_17__29_) );
  DFF_X2 decode_regfile_intregs_reg_17__30_ ( .D(n6740), .CK(clock), .Q(
        decode_regfile_intregs_17__30_) );
  DFF_X2 decode_regfile_intregs_reg_17__31_ ( .D(n6739), .CK(clock), .Q(
        decode_regfile_intregs_17__31_) );
  DFF_X2 decode_regfile_intregs_reg_16__0_ ( .D(n6738), .CK(clock), .Q(
        decode_regfile_intregs_16__0_) );
  DFF_X2 decode_regfile_intregs_reg_16__1_ ( .D(n6737), .CK(clock), .Q(
        decode_regfile_intregs_16__1_) );
  DFF_X2 decode_regfile_intregs_reg_16__2_ ( .D(n6736), .CK(clock), .Q(
        decode_regfile_intregs_16__2_) );
  DFF_X2 decode_regfile_intregs_reg_16__3_ ( .D(n6735), .CK(clock), .Q(
        decode_regfile_intregs_16__3_) );
  DFF_X2 decode_regfile_intregs_reg_16__4_ ( .D(n6734), .CK(clock), .Q(
        decode_regfile_intregs_16__4_) );
  DFF_X2 decode_regfile_intregs_reg_16__5_ ( .D(n6733), .CK(clock), .Q(
        decode_regfile_intregs_16__5_) );
  DFF_X2 decode_regfile_intregs_reg_16__6_ ( .D(n6732), .CK(clock), .Q(
        decode_regfile_intregs_16__6_) );
  DFF_X2 decode_regfile_intregs_reg_16__7_ ( .D(n6731), .CK(clock), .Q(
        decode_regfile_intregs_16__7_) );
  DFF_X2 decode_regfile_intregs_reg_16__8_ ( .D(n6730), .CK(clock), .Q(
        decode_regfile_intregs_16__8_) );
  DFF_X2 decode_regfile_intregs_reg_16__9_ ( .D(n6729), .CK(clock), .Q(
        decode_regfile_intregs_16__9_) );
  DFF_X2 decode_regfile_intregs_reg_16__10_ ( .D(n6728), .CK(clock), .Q(
        decode_regfile_intregs_16__10_) );
  DFF_X2 decode_regfile_intregs_reg_16__11_ ( .D(n6727), .CK(clock), .Q(
        decode_regfile_intregs_16__11_) );
  DFF_X2 decode_regfile_intregs_reg_16__12_ ( .D(n6726), .CK(clock), .Q(
        decode_regfile_intregs_16__12_) );
  DFF_X2 decode_regfile_intregs_reg_16__13_ ( .D(n6725), .CK(clock), .Q(
        decode_regfile_intregs_16__13_) );
  DFF_X2 decode_regfile_intregs_reg_16__14_ ( .D(n6724), .CK(clock), .Q(
        decode_regfile_intregs_16__14_) );
  DFF_X2 decode_regfile_intregs_reg_16__15_ ( .D(n6723), .CK(clock), .Q(
        decode_regfile_intregs_16__15_) );
  DFF_X2 decode_regfile_intregs_reg_16__16_ ( .D(n6722), .CK(clock), .Q(
        decode_regfile_intregs_16__16_) );
  DFF_X2 decode_regfile_intregs_reg_16__17_ ( .D(n6721), .CK(clock), .Q(
        decode_regfile_intregs_16__17_) );
  DFF_X2 decode_regfile_intregs_reg_16__18_ ( .D(n6720), .CK(clock), .Q(
        decode_regfile_intregs_16__18_) );
  DFF_X2 decode_regfile_intregs_reg_16__19_ ( .D(n6719), .CK(clock), .Q(
        decode_regfile_intregs_16__19_) );
  DFF_X2 decode_regfile_intregs_reg_16__20_ ( .D(n6718), .CK(clock), .Q(
        decode_regfile_intregs_16__20_) );
  DFF_X2 decode_regfile_intregs_reg_16__21_ ( .D(n6717), .CK(clock), .Q(
        decode_regfile_intregs_16__21_) );
  DFF_X2 decode_regfile_intregs_reg_16__22_ ( .D(n6716), .CK(clock), .Q(
        decode_regfile_intregs_16__22_) );
  DFF_X2 decode_regfile_intregs_reg_16__23_ ( .D(n6715), .CK(clock), .Q(
        decode_regfile_intregs_16__23_) );
  DFF_X2 decode_regfile_intregs_reg_16__24_ ( .D(n6714), .CK(clock), .Q(
        decode_regfile_intregs_16__24_) );
  DFF_X2 decode_regfile_intregs_reg_16__25_ ( .D(n6713), .CK(clock), .Q(
        decode_regfile_intregs_16__25_) );
  DFF_X2 decode_regfile_intregs_reg_16__26_ ( .D(n6712), .CK(clock), .Q(
        decode_regfile_intregs_16__26_) );
  DFF_X2 decode_regfile_intregs_reg_16__27_ ( .D(n6711), .CK(clock), .Q(
        decode_regfile_intregs_16__27_) );
  DFF_X2 decode_regfile_intregs_reg_16__28_ ( .D(n6710), .CK(clock), .Q(
        decode_regfile_intregs_16__28_) );
  DFF_X2 decode_regfile_intregs_reg_16__29_ ( .D(n6709), .CK(clock), .Q(
        decode_regfile_intregs_16__29_) );
  DFF_X2 decode_regfile_intregs_reg_16__30_ ( .D(n6708), .CK(clock), .Q(
        decode_regfile_intregs_16__30_) );
  DFF_X2 decode_regfile_intregs_reg_16__31_ ( .D(n6707), .CK(clock), .Q(
        decode_regfile_intregs_16__31_) );
  DFF_X2 decode_regfile_intregs_reg_15__0_ ( .D(n6706), .CK(clock), .Q(
        decode_regfile_intregs_15__0_) );
  DFF_X2 decode_regfile_intregs_reg_15__1_ ( .D(n6705), .CK(clock), .Q(
        decode_regfile_intregs_15__1_) );
  DFF_X2 decode_regfile_intregs_reg_15__2_ ( .D(n6704), .CK(clock), .Q(
        decode_regfile_intregs_15__2_) );
  DFF_X2 decode_regfile_intregs_reg_15__3_ ( .D(n6703), .CK(clock), .Q(
        decode_regfile_intregs_15__3_) );
  DFF_X2 decode_regfile_intregs_reg_15__4_ ( .D(n6702), .CK(clock), .Q(
        decode_regfile_intregs_15__4_) );
  DFF_X2 decode_regfile_intregs_reg_15__5_ ( .D(n6701), .CK(clock), .Q(
        decode_regfile_intregs_15__5_) );
  DFF_X2 decode_regfile_intregs_reg_15__6_ ( .D(n6700), .CK(clock), .Q(
        decode_regfile_intregs_15__6_) );
  DFF_X2 decode_regfile_intregs_reg_15__7_ ( .D(n6699), .CK(clock), .Q(
        decode_regfile_intregs_15__7_) );
  DFF_X2 decode_regfile_intregs_reg_15__8_ ( .D(n6698), .CK(clock), .Q(
        decode_regfile_intregs_15__8_) );
  DFF_X2 decode_regfile_intregs_reg_15__9_ ( .D(n6697), .CK(clock), .Q(
        decode_regfile_intregs_15__9_) );
  DFF_X2 decode_regfile_intregs_reg_15__10_ ( .D(n6696), .CK(clock), .Q(
        decode_regfile_intregs_15__10_) );
  DFF_X2 decode_regfile_intregs_reg_15__11_ ( .D(n6695), .CK(clock), .Q(
        decode_regfile_intregs_15__11_) );
  DFF_X2 decode_regfile_intregs_reg_15__12_ ( .D(n6694), .CK(clock), .Q(
        decode_regfile_intregs_15__12_) );
  DFF_X2 decode_regfile_intregs_reg_15__13_ ( .D(n6693), .CK(clock), .Q(
        decode_regfile_intregs_15__13_) );
  DFF_X2 decode_regfile_intregs_reg_15__14_ ( .D(n6692), .CK(clock), .Q(
        decode_regfile_intregs_15__14_) );
  DFF_X2 decode_regfile_intregs_reg_15__15_ ( .D(n6691), .CK(clock), .Q(
        decode_regfile_intregs_15__15_) );
  DFF_X2 decode_regfile_intregs_reg_15__16_ ( .D(n6690), .CK(clock), .Q(
        decode_regfile_intregs_15__16_) );
  DFF_X2 decode_regfile_intregs_reg_15__17_ ( .D(n6689), .CK(clock), .Q(
        decode_regfile_intregs_15__17_) );
  DFF_X2 decode_regfile_intregs_reg_15__18_ ( .D(n6688), .CK(clock), .Q(
        decode_regfile_intregs_15__18_) );
  DFF_X2 decode_regfile_intregs_reg_15__19_ ( .D(n6687), .CK(clock), .Q(
        decode_regfile_intregs_15__19_) );
  DFF_X2 decode_regfile_intregs_reg_15__20_ ( .D(n6686), .CK(clock), .Q(
        decode_regfile_intregs_15__20_) );
  DFF_X2 decode_regfile_intregs_reg_15__21_ ( .D(n6685), .CK(clock), .Q(
        decode_regfile_intregs_15__21_) );
  DFF_X2 decode_regfile_intregs_reg_15__22_ ( .D(n6684), .CK(clock), .Q(
        decode_regfile_intregs_15__22_) );
  DFF_X2 decode_regfile_intregs_reg_15__23_ ( .D(n6683), .CK(clock), .Q(
        decode_regfile_intregs_15__23_) );
  DFF_X2 decode_regfile_intregs_reg_15__24_ ( .D(n6682), .CK(clock), .Q(
        decode_regfile_intregs_15__24_) );
  DFF_X2 decode_regfile_intregs_reg_15__25_ ( .D(n6681), .CK(clock), .Q(
        decode_regfile_intregs_15__25_) );
  DFF_X2 decode_regfile_intregs_reg_15__26_ ( .D(n6680), .CK(clock), .Q(
        decode_regfile_intregs_15__26_) );
  DFF_X2 decode_regfile_intregs_reg_15__27_ ( .D(n6679), .CK(clock), .Q(
        decode_regfile_intregs_15__27_) );
  DFF_X2 decode_regfile_intregs_reg_15__28_ ( .D(n6678), .CK(clock), .Q(
        decode_regfile_intregs_15__28_) );
  DFF_X2 decode_regfile_intregs_reg_15__29_ ( .D(n6677), .CK(clock), .Q(
        decode_regfile_intregs_15__29_) );
  DFF_X2 decode_regfile_intregs_reg_15__30_ ( .D(n6676), .CK(clock), .Q(
        decode_regfile_intregs_15__30_) );
  DFF_X2 decode_regfile_intregs_reg_15__31_ ( .D(n6675), .CK(clock), .Q(
        decode_regfile_intregs_15__31_) );
  DFF_X2 decode_regfile_intregs_reg_14__0_ ( .D(n6674), .CK(clock), .Q(
        decode_regfile_intregs_14__0_) );
  DFF_X2 decode_regfile_intregs_reg_14__1_ ( .D(n6673), .CK(clock), .Q(
        decode_regfile_intregs_14__1_) );
  DFF_X2 decode_regfile_intregs_reg_14__2_ ( .D(n6672), .CK(clock), .Q(
        decode_regfile_intregs_14__2_) );
  DFF_X2 decode_regfile_intregs_reg_14__3_ ( .D(n6671), .CK(clock), .Q(
        decode_regfile_intregs_14__3_) );
  DFF_X2 decode_regfile_intregs_reg_14__4_ ( .D(n6670), .CK(clock), .Q(
        decode_regfile_intregs_14__4_) );
  DFF_X2 decode_regfile_intregs_reg_14__5_ ( .D(n6669), .CK(clock), .Q(
        decode_regfile_intregs_14__5_) );
  DFF_X2 decode_regfile_intregs_reg_14__6_ ( .D(n6668), .CK(clock), .Q(
        decode_regfile_intregs_14__6_) );
  DFF_X2 decode_regfile_intregs_reg_14__7_ ( .D(n6667), .CK(clock), .Q(
        decode_regfile_intregs_14__7_) );
  DFF_X2 decode_regfile_intregs_reg_14__8_ ( .D(n6666), .CK(clock), .Q(
        decode_regfile_intregs_14__8_) );
  DFF_X2 decode_regfile_intregs_reg_14__9_ ( .D(n6665), .CK(clock), .Q(
        decode_regfile_intregs_14__9_) );
  DFF_X2 decode_regfile_intregs_reg_14__10_ ( .D(n6664), .CK(clock), .Q(
        decode_regfile_intregs_14__10_) );
  DFF_X2 decode_regfile_intregs_reg_14__11_ ( .D(n6663), .CK(clock), .Q(
        decode_regfile_intregs_14__11_) );
  DFF_X2 decode_regfile_intregs_reg_14__12_ ( .D(n6662), .CK(clock), .Q(
        decode_regfile_intregs_14__12_) );
  DFF_X2 decode_regfile_intregs_reg_14__13_ ( .D(n6661), .CK(clock), .Q(
        decode_regfile_intregs_14__13_) );
  DFF_X2 decode_regfile_intregs_reg_14__14_ ( .D(n6660), .CK(clock), .Q(
        decode_regfile_intregs_14__14_) );
  DFF_X2 decode_regfile_intregs_reg_14__15_ ( .D(n6659), .CK(clock), .Q(
        decode_regfile_intregs_14__15_) );
  DFF_X2 decode_regfile_intregs_reg_14__16_ ( .D(n6658), .CK(clock), .Q(
        decode_regfile_intregs_14__16_) );
  DFF_X2 decode_regfile_intregs_reg_14__17_ ( .D(n6657), .CK(clock), .Q(
        decode_regfile_intregs_14__17_) );
  DFF_X2 decode_regfile_intregs_reg_14__18_ ( .D(n6656), .CK(clock), .Q(
        decode_regfile_intregs_14__18_) );
  DFF_X2 decode_regfile_intregs_reg_14__19_ ( .D(n6655), .CK(clock), .Q(
        decode_regfile_intregs_14__19_) );
  DFF_X2 decode_regfile_intregs_reg_14__20_ ( .D(n6654), .CK(clock), .Q(
        decode_regfile_intregs_14__20_) );
  DFF_X2 decode_regfile_intregs_reg_14__21_ ( .D(n6653), .CK(clock), .Q(
        decode_regfile_intregs_14__21_) );
  DFF_X2 decode_regfile_intregs_reg_14__22_ ( .D(n6652), .CK(clock), .Q(
        decode_regfile_intregs_14__22_) );
  DFF_X2 decode_regfile_intregs_reg_14__23_ ( .D(n6651), .CK(clock), .Q(
        decode_regfile_intregs_14__23_) );
  DFF_X2 decode_regfile_intregs_reg_14__24_ ( .D(n6650), .CK(clock), .Q(
        decode_regfile_intregs_14__24_) );
  DFF_X2 decode_regfile_intregs_reg_14__25_ ( .D(n6649), .CK(clock), .Q(
        decode_regfile_intregs_14__25_) );
  DFF_X2 decode_regfile_intregs_reg_14__26_ ( .D(n6648), .CK(clock), .Q(
        decode_regfile_intregs_14__26_) );
  DFF_X2 decode_regfile_intregs_reg_14__27_ ( .D(n6647), .CK(clock), .Q(
        decode_regfile_intregs_14__27_) );
  DFF_X2 decode_regfile_intregs_reg_14__28_ ( .D(n6646), .CK(clock), .Q(
        decode_regfile_intregs_14__28_) );
  DFF_X2 decode_regfile_intregs_reg_14__29_ ( .D(n6645), .CK(clock), .Q(
        decode_regfile_intregs_14__29_) );
  DFF_X2 decode_regfile_intregs_reg_14__30_ ( .D(n6644), .CK(clock), .Q(
        decode_regfile_intregs_14__30_) );
  DFF_X2 decode_regfile_intregs_reg_14__31_ ( .D(n6643), .CK(clock), .Q(
        decode_regfile_intregs_14__31_) );
  DFF_X2 decode_regfile_intregs_reg_13__0_ ( .D(n6642), .CK(clock), .Q(
        decode_regfile_intregs_13__0_) );
  DFF_X2 decode_regfile_intregs_reg_13__1_ ( .D(n6641), .CK(clock), .Q(
        decode_regfile_intregs_13__1_) );
  DFF_X2 decode_regfile_intregs_reg_13__2_ ( .D(n6640), .CK(clock), .Q(
        decode_regfile_intregs_13__2_) );
  DFF_X2 decode_regfile_intregs_reg_13__3_ ( .D(n6639), .CK(clock), .Q(
        decode_regfile_intregs_13__3_) );
  DFF_X2 decode_regfile_intregs_reg_13__4_ ( .D(n6638), .CK(clock), .Q(
        decode_regfile_intregs_13__4_) );
  DFF_X2 decode_regfile_intregs_reg_13__5_ ( .D(n6637), .CK(clock), .Q(
        decode_regfile_intregs_13__5_) );
  DFF_X2 decode_regfile_intregs_reg_13__6_ ( .D(n6636), .CK(clock), .Q(
        decode_regfile_intregs_13__6_) );
  DFF_X2 decode_regfile_intregs_reg_13__7_ ( .D(n6635), .CK(clock), .Q(
        decode_regfile_intregs_13__7_) );
  DFF_X2 decode_regfile_intregs_reg_13__8_ ( .D(n6634), .CK(clock), .Q(
        decode_regfile_intregs_13__8_) );
  DFF_X2 decode_regfile_intregs_reg_13__9_ ( .D(n6633), .CK(clock), .Q(
        decode_regfile_intregs_13__9_) );
  DFF_X2 decode_regfile_intregs_reg_13__10_ ( .D(n6632), .CK(clock), .Q(
        decode_regfile_intregs_13__10_) );
  DFF_X2 decode_regfile_intregs_reg_13__11_ ( .D(n6631), .CK(clock), .Q(
        decode_regfile_intregs_13__11_) );
  DFF_X2 decode_regfile_intregs_reg_13__12_ ( .D(n6630), .CK(clock), .Q(
        decode_regfile_intregs_13__12_) );
  DFF_X2 decode_regfile_intregs_reg_13__13_ ( .D(n6629), .CK(clock), .Q(
        decode_regfile_intregs_13__13_) );
  DFF_X2 decode_regfile_intregs_reg_13__14_ ( .D(n6628), .CK(clock), .Q(
        decode_regfile_intregs_13__14_) );
  DFF_X2 decode_regfile_intregs_reg_13__15_ ( .D(n6627), .CK(clock), .Q(
        decode_regfile_intregs_13__15_) );
  DFF_X2 decode_regfile_intregs_reg_13__16_ ( .D(n6626), .CK(clock), .Q(
        decode_regfile_intregs_13__16_) );
  DFF_X2 decode_regfile_intregs_reg_13__17_ ( .D(n6625), .CK(clock), .Q(
        decode_regfile_intregs_13__17_) );
  DFF_X2 decode_regfile_intregs_reg_13__18_ ( .D(n6624), .CK(clock), .Q(
        decode_regfile_intregs_13__18_) );
  DFF_X2 decode_regfile_intregs_reg_13__19_ ( .D(n6623), .CK(clock), .Q(
        decode_regfile_intregs_13__19_) );
  DFF_X2 decode_regfile_intregs_reg_13__20_ ( .D(n6622), .CK(clock), .Q(
        decode_regfile_intregs_13__20_) );
  DFF_X2 decode_regfile_intregs_reg_13__21_ ( .D(n6621), .CK(clock), .Q(
        decode_regfile_intregs_13__21_) );
  DFF_X2 decode_regfile_intregs_reg_13__22_ ( .D(n6620), .CK(clock), .Q(
        decode_regfile_intregs_13__22_) );
  DFF_X2 decode_regfile_intregs_reg_13__23_ ( .D(n6619), .CK(clock), .Q(
        decode_regfile_intregs_13__23_) );
  DFF_X2 decode_regfile_intregs_reg_13__24_ ( .D(n6618), .CK(clock), .Q(
        decode_regfile_intregs_13__24_) );
  DFF_X2 decode_regfile_intregs_reg_13__25_ ( .D(n6617), .CK(clock), .Q(
        decode_regfile_intregs_13__25_) );
  DFF_X2 decode_regfile_intregs_reg_13__26_ ( .D(n6616), .CK(clock), .Q(
        decode_regfile_intregs_13__26_) );
  DFF_X2 decode_regfile_intregs_reg_13__27_ ( .D(n6615), .CK(clock), .Q(
        decode_regfile_intregs_13__27_) );
  DFF_X2 decode_regfile_intregs_reg_13__28_ ( .D(n6614), .CK(clock), .Q(
        decode_regfile_intregs_13__28_) );
  DFF_X2 decode_regfile_intregs_reg_13__29_ ( .D(n6613), .CK(clock), .Q(
        decode_regfile_intregs_13__29_) );
  DFF_X2 decode_regfile_intregs_reg_13__30_ ( .D(n6612), .CK(clock), .Q(
        decode_regfile_intregs_13__30_) );
  DFF_X2 decode_regfile_intregs_reg_13__31_ ( .D(n6611), .CK(clock), .Q(
        decode_regfile_intregs_13__31_) );
  DFF_X2 decode_regfile_intregs_reg_12__0_ ( .D(n6610), .CK(clock), .Q(
        decode_regfile_intregs_12__0_) );
  DFF_X2 decode_regfile_intregs_reg_12__1_ ( .D(n6609), .CK(clock), .Q(
        decode_regfile_intregs_12__1_) );
  DFF_X2 decode_regfile_intregs_reg_12__2_ ( .D(n6608), .CK(clock), .Q(
        decode_regfile_intregs_12__2_) );
  DFF_X2 decode_regfile_intregs_reg_12__3_ ( .D(n6607), .CK(clock), .Q(
        decode_regfile_intregs_12__3_) );
  DFF_X2 decode_regfile_intregs_reg_12__4_ ( .D(n6606), .CK(clock), .Q(
        decode_regfile_intregs_12__4_) );
  DFF_X2 decode_regfile_intregs_reg_12__5_ ( .D(n6605), .CK(clock), .Q(
        decode_regfile_intregs_12__5_) );
  DFF_X2 decode_regfile_intregs_reg_12__6_ ( .D(n6604), .CK(clock), .Q(
        decode_regfile_intregs_12__6_) );
  DFF_X2 decode_regfile_intregs_reg_12__7_ ( .D(n6603), .CK(clock), .Q(
        decode_regfile_intregs_12__7_) );
  DFF_X2 decode_regfile_intregs_reg_12__8_ ( .D(n6602), .CK(clock), .Q(
        decode_regfile_intregs_12__8_) );
  DFF_X2 decode_regfile_intregs_reg_12__9_ ( .D(n6601), .CK(clock), .Q(
        decode_regfile_intregs_12__9_) );
  DFF_X2 decode_regfile_intregs_reg_12__10_ ( .D(n6600), .CK(clock), .Q(
        decode_regfile_intregs_12__10_) );
  DFF_X2 decode_regfile_intregs_reg_12__11_ ( .D(n6599), .CK(clock), .Q(
        decode_regfile_intregs_12__11_) );
  DFF_X2 decode_regfile_intregs_reg_12__12_ ( .D(n6598), .CK(clock), .Q(
        decode_regfile_intregs_12__12_) );
  DFF_X2 decode_regfile_intregs_reg_12__13_ ( .D(n6597), .CK(clock), .Q(
        decode_regfile_intregs_12__13_) );
  DFF_X2 decode_regfile_intregs_reg_12__14_ ( .D(n6596), .CK(clock), .Q(
        decode_regfile_intregs_12__14_) );
  DFF_X2 decode_regfile_intregs_reg_12__15_ ( .D(n6595), .CK(clock), .Q(
        decode_regfile_intregs_12__15_) );
  DFF_X2 decode_regfile_intregs_reg_12__16_ ( .D(n6594), .CK(clock), .Q(
        decode_regfile_intregs_12__16_) );
  DFF_X2 decode_regfile_intregs_reg_12__17_ ( .D(n6593), .CK(clock), .Q(
        decode_regfile_intregs_12__17_) );
  DFF_X2 decode_regfile_intregs_reg_12__18_ ( .D(n6592), .CK(clock), .Q(
        decode_regfile_intregs_12__18_) );
  DFF_X2 decode_regfile_intregs_reg_12__19_ ( .D(n6591), .CK(clock), .Q(
        decode_regfile_intregs_12__19_) );
  DFF_X2 decode_regfile_intregs_reg_12__20_ ( .D(n6590), .CK(clock), .Q(
        decode_regfile_intregs_12__20_) );
  DFF_X2 decode_regfile_intregs_reg_12__21_ ( .D(n6589), .CK(clock), .Q(
        decode_regfile_intregs_12__21_) );
  DFF_X2 decode_regfile_intregs_reg_12__22_ ( .D(n6588), .CK(clock), .Q(
        decode_regfile_intregs_12__22_) );
  DFF_X2 decode_regfile_intregs_reg_12__23_ ( .D(n6587), .CK(clock), .Q(
        decode_regfile_intregs_12__23_) );
  DFF_X2 decode_regfile_intregs_reg_12__24_ ( .D(n6586), .CK(clock), .Q(
        decode_regfile_intregs_12__24_) );
  DFF_X2 decode_regfile_intregs_reg_12__25_ ( .D(n6585), .CK(clock), .Q(
        decode_regfile_intregs_12__25_) );
  DFF_X2 decode_regfile_intregs_reg_12__26_ ( .D(n6584), .CK(clock), .Q(
        decode_regfile_intregs_12__26_) );
  DFF_X2 decode_regfile_intregs_reg_12__27_ ( .D(n6583), .CK(clock), .Q(
        decode_regfile_intregs_12__27_) );
  DFF_X2 decode_regfile_intregs_reg_12__28_ ( .D(n6582), .CK(clock), .Q(
        decode_regfile_intregs_12__28_) );
  DFF_X2 decode_regfile_intregs_reg_12__29_ ( .D(n6581), .CK(clock), .Q(
        decode_regfile_intregs_12__29_) );
  DFF_X2 decode_regfile_intregs_reg_12__30_ ( .D(n6580), .CK(clock), .Q(
        decode_regfile_intregs_12__30_) );
  DFF_X2 decode_regfile_intregs_reg_12__31_ ( .D(n6579), .CK(clock), .Q(
        decode_regfile_intregs_12__31_) );
  DFF_X2 decode_regfile_intregs_reg_11__0_ ( .D(n6578), .CK(clock), .Q(
        decode_regfile_intregs_11__0_) );
  DFF_X2 decode_regfile_intregs_reg_11__1_ ( .D(n6577), .CK(clock), .Q(
        decode_regfile_intregs_11__1_) );
  DFF_X2 decode_regfile_intregs_reg_11__2_ ( .D(n6576), .CK(clock), .Q(
        decode_regfile_intregs_11__2_) );
  DFF_X2 decode_regfile_intregs_reg_11__3_ ( .D(n6575), .CK(clock), .Q(
        decode_regfile_intregs_11__3_) );
  DFF_X2 decode_regfile_intregs_reg_11__4_ ( .D(n6574), .CK(clock), .Q(
        decode_regfile_intregs_11__4_) );
  DFF_X2 decode_regfile_intregs_reg_11__5_ ( .D(n6573), .CK(clock), .Q(
        decode_regfile_intregs_11__5_) );
  DFF_X2 decode_regfile_intregs_reg_11__6_ ( .D(n6572), .CK(clock), .Q(
        decode_regfile_intregs_11__6_) );
  DFF_X2 decode_regfile_intregs_reg_11__7_ ( .D(n6571), .CK(clock), .Q(
        decode_regfile_intregs_11__7_) );
  DFF_X2 decode_regfile_intregs_reg_11__8_ ( .D(n6570), .CK(clock), .Q(
        decode_regfile_intregs_11__8_) );
  DFF_X2 decode_regfile_intregs_reg_11__9_ ( .D(n6569), .CK(clock), .Q(
        decode_regfile_intregs_11__9_) );
  DFF_X2 decode_regfile_intregs_reg_11__10_ ( .D(n6568), .CK(clock), .Q(
        decode_regfile_intregs_11__10_) );
  DFF_X2 decode_regfile_intregs_reg_11__11_ ( .D(n6567), .CK(clock), .Q(
        decode_regfile_intregs_11__11_) );
  DFF_X2 decode_regfile_intregs_reg_11__12_ ( .D(n6566), .CK(clock), .Q(
        decode_regfile_intregs_11__12_) );
  DFF_X2 decode_regfile_intregs_reg_11__13_ ( .D(n6565), .CK(clock), .Q(
        decode_regfile_intregs_11__13_) );
  DFF_X2 decode_regfile_intregs_reg_11__14_ ( .D(n6564), .CK(clock), .Q(
        decode_regfile_intregs_11__14_) );
  DFF_X2 decode_regfile_intregs_reg_11__15_ ( .D(n6563), .CK(clock), .Q(
        decode_regfile_intregs_11__15_) );
  DFF_X2 decode_regfile_intregs_reg_11__16_ ( .D(n6562), .CK(clock), .Q(
        decode_regfile_intregs_11__16_) );
  DFF_X2 decode_regfile_intregs_reg_11__17_ ( .D(n6561), .CK(clock), .Q(
        decode_regfile_intregs_11__17_) );
  DFF_X2 decode_regfile_intregs_reg_11__18_ ( .D(n6560), .CK(clock), .Q(
        decode_regfile_intregs_11__18_) );
  DFF_X2 decode_regfile_intregs_reg_11__19_ ( .D(n6559), .CK(clock), .Q(
        decode_regfile_intregs_11__19_) );
  DFF_X2 decode_regfile_intregs_reg_11__20_ ( .D(n6558), .CK(clock), .Q(
        decode_regfile_intregs_11__20_) );
  DFF_X2 decode_regfile_intregs_reg_11__21_ ( .D(n6557), .CK(clock), .Q(
        decode_regfile_intregs_11__21_) );
  DFF_X2 decode_regfile_intregs_reg_11__22_ ( .D(n6556), .CK(clock), .Q(
        decode_regfile_intregs_11__22_) );
  DFF_X2 decode_regfile_intregs_reg_11__23_ ( .D(n6555), .CK(clock), .Q(
        decode_regfile_intregs_11__23_) );
  DFF_X2 decode_regfile_intregs_reg_11__24_ ( .D(n6554), .CK(clock), .Q(
        decode_regfile_intregs_11__24_) );
  DFF_X2 decode_regfile_intregs_reg_11__25_ ( .D(n6553), .CK(clock), .Q(
        decode_regfile_intregs_11__25_) );
  DFF_X2 decode_regfile_intregs_reg_11__26_ ( .D(n6552), .CK(clock), .Q(
        decode_regfile_intregs_11__26_) );
  DFF_X2 decode_regfile_intregs_reg_11__27_ ( .D(n6551), .CK(clock), .Q(
        decode_regfile_intregs_11__27_) );
  DFF_X2 decode_regfile_intregs_reg_11__28_ ( .D(n6550), .CK(clock), .Q(
        decode_regfile_intregs_11__28_) );
  DFF_X2 decode_regfile_intregs_reg_11__29_ ( .D(n6549), .CK(clock), .Q(
        decode_regfile_intregs_11__29_) );
  DFF_X2 decode_regfile_intregs_reg_11__30_ ( .D(n6548), .CK(clock), .Q(
        decode_regfile_intregs_11__30_) );
  DFF_X2 decode_regfile_intregs_reg_11__31_ ( .D(n6547), .CK(clock), .Q(
        decode_regfile_intregs_11__31_) );
  DFF_X2 decode_regfile_intregs_reg_10__0_ ( .D(n6546), .CK(clock), .Q(
        decode_regfile_intregs_10__0_) );
  DFF_X2 decode_regfile_intregs_reg_10__1_ ( .D(n6545), .CK(clock), .Q(
        decode_regfile_intregs_10__1_) );
  DFF_X2 decode_regfile_intregs_reg_10__2_ ( .D(n6544), .CK(clock), .Q(
        decode_regfile_intregs_10__2_) );
  DFF_X2 decode_regfile_intregs_reg_10__3_ ( .D(n6543), .CK(clock), .Q(
        decode_regfile_intregs_10__3_) );
  DFF_X2 decode_regfile_intregs_reg_10__4_ ( .D(n6542), .CK(clock), .Q(
        decode_regfile_intregs_10__4_) );
  DFF_X2 decode_regfile_intregs_reg_10__5_ ( .D(n6541), .CK(clock), .Q(
        decode_regfile_intregs_10__5_) );
  DFF_X2 decode_regfile_intregs_reg_10__6_ ( .D(n6540), .CK(clock), .Q(
        decode_regfile_intregs_10__6_) );
  DFF_X2 decode_regfile_intregs_reg_10__7_ ( .D(n6539), .CK(clock), .Q(
        decode_regfile_intregs_10__7_) );
  DFF_X2 decode_regfile_intregs_reg_10__8_ ( .D(n6538), .CK(clock), .Q(
        decode_regfile_intregs_10__8_) );
  DFF_X2 decode_regfile_intregs_reg_10__9_ ( .D(n6537), .CK(clock), .Q(
        decode_regfile_intregs_10__9_) );
  DFF_X2 decode_regfile_intregs_reg_10__10_ ( .D(n6536), .CK(clock), .Q(
        decode_regfile_intregs_10__10_) );
  DFF_X2 decode_regfile_intregs_reg_10__11_ ( .D(n6535), .CK(clock), .Q(
        decode_regfile_intregs_10__11_) );
  DFF_X2 decode_regfile_intregs_reg_10__12_ ( .D(n6534), .CK(clock), .Q(
        decode_regfile_intregs_10__12_) );
  DFF_X2 decode_regfile_intregs_reg_10__13_ ( .D(n6533), .CK(clock), .Q(
        decode_regfile_intregs_10__13_) );
  DFF_X2 decode_regfile_intregs_reg_10__14_ ( .D(n6532), .CK(clock), .Q(
        decode_regfile_intregs_10__14_) );
  DFF_X2 decode_regfile_intregs_reg_10__15_ ( .D(n6531), .CK(clock), .Q(
        decode_regfile_intregs_10__15_) );
  DFF_X2 decode_regfile_intregs_reg_10__16_ ( .D(n6530), .CK(clock), .Q(
        decode_regfile_intregs_10__16_) );
  DFF_X2 decode_regfile_intregs_reg_10__17_ ( .D(n6529), .CK(clock), .Q(
        decode_regfile_intregs_10__17_) );
  DFF_X2 decode_regfile_intregs_reg_10__18_ ( .D(n6528), .CK(clock), .Q(
        decode_regfile_intregs_10__18_) );
  DFF_X2 decode_regfile_intregs_reg_10__19_ ( .D(n6527), .CK(clock), .Q(
        decode_regfile_intregs_10__19_) );
  DFF_X2 decode_regfile_intregs_reg_10__20_ ( .D(n6526), .CK(clock), .Q(
        decode_regfile_intregs_10__20_) );
  DFF_X2 decode_regfile_intregs_reg_10__21_ ( .D(n6525), .CK(clock), .Q(
        decode_regfile_intregs_10__21_) );
  DFF_X2 decode_regfile_intregs_reg_10__22_ ( .D(n6524), .CK(clock), .Q(
        decode_regfile_intregs_10__22_) );
  DFF_X2 decode_regfile_intregs_reg_10__23_ ( .D(n6523), .CK(clock), .Q(
        decode_regfile_intregs_10__23_) );
  DFF_X2 decode_regfile_intregs_reg_10__24_ ( .D(n6522), .CK(clock), .Q(
        decode_regfile_intregs_10__24_) );
  DFF_X2 decode_regfile_intregs_reg_10__25_ ( .D(n6521), .CK(clock), .Q(
        decode_regfile_intregs_10__25_) );
  DFF_X2 decode_regfile_intregs_reg_10__26_ ( .D(n6520), .CK(clock), .Q(
        decode_regfile_intregs_10__26_) );
  DFF_X2 decode_regfile_intregs_reg_10__27_ ( .D(n6519), .CK(clock), .Q(
        decode_regfile_intregs_10__27_) );
  DFF_X2 decode_regfile_intregs_reg_10__28_ ( .D(n6518), .CK(clock), .Q(
        decode_regfile_intregs_10__28_) );
  DFF_X2 decode_regfile_intregs_reg_10__29_ ( .D(n6517), .CK(clock), .Q(
        decode_regfile_intregs_10__29_) );
  DFF_X2 decode_regfile_intregs_reg_10__30_ ( .D(n6516), .CK(clock), .Q(
        decode_regfile_intregs_10__30_) );
  DFF_X2 decode_regfile_intregs_reg_10__31_ ( .D(n6515), .CK(clock), .Q(
        decode_regfile_intregs_10__31_) );
  DFF_X2 decode_regfile_intregs_reg_9__0_ ( .D(n6514), .CK(clock), .Q(
        decode_regfile_intregs_9__0_) );
  DFF_X2 decode_regfile_intregs_reg_9__1_ ( .D(n6513), .CK(clock), .Q(
        decode_regfile_intregs_9__1_) );
  DFF_X2 decode_regfile_intregs_reg_9__2_ ( .D(n6512), .CK(clock), .Q(
        decode_regfile_intregs_9__2_) );
  DFF_X2 decode_regfile_intregs_reg_9__3_ ( .D(n6511), .CK(clock), .Q(
        decode_regfile_intregs_9__3_) );
  DFF_X2 decode_regfile_intregs_reg_9__4_ ( .D(n6510), .CK(clock), .Q(
        decode_regfile_intregs_9__4_) );
  DFF_X2 decode_regfile_intregs_reg_9__5_ ( .D(n6509), .CK(clock), .Q(
        decode_regfile_intregs_9__5_) );
  DFF_X2 decode_regfile_intregs_reg_9__6_ ( .D(n6508), .CK(clock), .Q(
        decode_regfile_intregs_9__6_) );
  DFF_X2 decode_regfile_intregs_reg_9__7_ ( .D(n6507), .CK(clock), .Q(
        decode_regfile_intregs_9__7_) );
  DFF_X2 decode_regfile_intregs_reg_9__8_ ( .D(n6506), .CK(clock), .Q(
        decode_regfile_intregs_9__8_) );
  DFF_X2 decode_regfile_intregs_reg_9__9_ ( .D(n6505), .CK(clock), .Q(
        decode_regfile_intregs_9__9_) );
  DFF_X2 decode_regfile_intregs_reg_9__10_ ( .D(n6504), .CK(clock), .Q(
        decode_regfile_intregs_9__10_) );
  DFF_X2 decode_regfile_intregs_reg_9__11_ ( .D(n6503), .CK(clock), .Q(
        decode_regfile_intregs_9__11_) );
  DFF_X2 decode_regfile_intregs_reg_9__12_ ( .D(n6502), .CK(clock), .Q(
        decode_regfile_intregs_9__12_) );
  DFF_X2 decode_regfile_intregs_reg_9__13_ ( .D(n6501), .CK(clock), .Q(
        decode_regfile_intregs_9__13_) );
  DFF_X2 decode_regfile_intregs_reg_9__14_ ( .D(n6500), .CK(clock), .Q(
        decode_regfile_intregs_9__14_) );
  DFF_X2 decode_regfile_intregs_reg_9__15_ ( .D(n6499), .CK(clock), .Q(
        decode_regfile_intregs_9__15_) );
  DFF_X2 decode_regfile_intregs_reg_9__16_ ( .D(n6498), .CK(clock), .Q(
        decode_regfile_intregs_9__16_) );
  DFF_X2 decode_regfile_intregs_reg_9__17_ ( .D(n6497), .CK(clock), .Q(
        decode_regfile_intregs_9__17_) );
  DFF_X2 decode_regfile_intregs_reg_9__18_ ( .D(n6496), .CK(clock), .Q(
        decode_regfile_intregs_9__18_) );
  DFF_X2 decode_regfile_intregs_reg_9__19_ ( .D(n6495), .CK(clock), .Q(
        decode_regfile_intregs_9__19_) );
  DFF_X2 decode_regfile_intregs_reg_9__20_ ( .D(n6494), .CK(clock), .Q(
        decode_regfile_intregs_9__20_) );
  DFF_X2 decode_regfile_intregs_reg_9__21_ ( .D(n6493), .CK(clock), .Q(
        decode_regfile_intregs_9__21_) );
  DFF_X2 decode_regfile_intregs_reg_9__22_ ( .D(n6492), .CK(clock), .Q(
        decode_regfile_intregs_9__22_) );
  DFF_X2 decode_regfile_intregs_reg_9__23_ ( .D(n6491), .CK(clock), .Q(
        decode_regfile_intregs_9__23_) );
  DFF_X2 decode_regfile_intregs_reg_9__24_ ( .D(n6490), .CK(clock), .Q(
        decode_regfile_intregs_9__24_) );
  DFF_X2 decode_regfile_intregs_reg_9__25_ ( .D(n6489), .CK(clock), .Q(
        decode_regfile_intregs_9__25_) );
  DFF_X2 decode_regfile_intregs_reg_9__26_ ( .D(n6488), .CK(clock), .Q(
        decode_regfile_intregs_9__26_) );
  DFF_X2 decode_regfile_intregs_reg_9__27_ ( .D(n6487), .CK(clock), .Q(
        decode_regfile_intregs_9__27_) );
  DFF_X2 decode_regfile_intregs_reg_9__28_ ( .D(n6486), .CK(clock), .Q(
        decode_regfile_intregs_9__28_) );
  DFF_X2 decode_regfile_intregs_reg_9__29_ ( .D(n6485), .CK(clock), .Q(
        decode_regfile_intregs_9__29_) );
  DFF_X2 decode_regfile_intregs_reg_9__30_ ( .D(n6484), .CK(clock), .Q(
        decode_regfile_intregs_9__30_) );
  DFF_X2 decode_regfile_intregs_reg_9__31_ ( .D(n6483), .CK(clock), .Q(
        decode_regfile_intregs_9__31_) );
  DFF_X2 decode_regfile_intregs_reg_8__0_ ( .D(n6482), .CK(clock), .Q(
        decode_regfile_intregs_8__0_) );
  DFF_X2 decode_regfile_intregs_reg_8__1_ ( .D(n6481), .CK(clock), .Q(
        decode_regfile_intregs_8__1_) );
  DFF_X2 decode_regfile_intregs_reg_8__2_ ( .D(n6480), .CK(clock), .Q(
        decode_regfile_intregs_8__2_) );
  DFF_X2 decode_regfile_intregs_reg_8__3_ ( .D(n6479), .CK(clock), .Q(
        decode_regfile_intregs_8__3_) );
  DFF_X2 decode_regfile_intregs_reg_8__4_ ( .D(n6478), .CK(clock), .Q(
        decode_regfile_intregs_8__4_) );
  DFF_X2 decode_regfile_intregs_reg_8__5_ ( .D(n6477), .CK(clock), .Q(
        decode_regfile_intregs_8__5_) );
  DFF_X2 decode_regfile_intregs_reg_8__6_ ( .D(n6476), .CK(clock), .Q(
        decode_regfile_intregs_8__6_) );
  DFF_X2 decode_regfile_intregs_reg_8__7_ ( .D(n6475), .CK(clock), .Q(
        decode_regfile_intregs_8__7_) );
  DFF_X2 decode_regfile_intregs_reg_8__8_ ( .D(n6474), .CK(clock), .Q(
        decode_regfile_intregs_8__8_) );
  DFF_X2 decode_regfile_intregs_reg_8__9_ ( .D(n6473), .CK(clock), .Q(
        decode_regfile_intregs_8__9_) );
  DFF_X2 decode_regfile_intregs_reg_8__10_ ( .D(n6472), .CK(clock), .Q(
        decode_regfile_intregs_8__10_) );
  DFF_X2 decode_regfile_intregs_reg_8__11_ ( .D(n6471), .CK(clock), .Q(
        decode_regfile_intregs_8__11_) );
  DFF_X2 decode_regfile_intregs_reg_8__12_ ( .D(n6470), .CK(clock), .Q(
        decode_regfile_intregs_8__12_) );
  DFF_X2 decode_regfile_intregs_reg_8__13_ ( .D(n6469), .CK(clock), .Q(
        decode_regfile_intregs_8__13_) );
  DFF_X2 decode_regfile_intregs_reg_8__14_ ( .D(n6468), .CK(clock), .Q(
        decode_regfile_intregs_8__14_) );
  DFF_X2 decode_regfile_intregs_reg_8__15_ ( .D(n6467), .CK(clock), .Q(
        decode_regfile_intregs_8__15_) );
  DFF_X2 decode_regfile_intregs_reg_8__16_ ( .D(n6466), .CK(clock), .Q(
        decode_regfile_intregs_8__16_) );
  DFF_X2 decode_regfile_intregs_reg_8__17_ ( .D(n6465), .CK(clock), .Q(
        decode_regfile_intregs_8__17_) );
  DFF_X2 decode_regfile_intregs_reg_8__18_ ( .D(n6464), .CK(clock), .Q(
        decode_regfile_intregs_8__18_) );
  DFF_X2 decode_regfile_intregs_reg_8__19_ ( .D(n6463), .CK(clock), .Q(
        decode_regfile_intregs_8__19_) );
  DFF_X2 decode_regfile_intregs_reg_8__20_ ( .D(n6462), .CK(clock), .Q(
        decode_regfile_intregs_8__20_) );
  DFF_X2 decode_regfile_intregs_reg_8__21_ ( .D(n6461), .CK(clock), .Q(
        decode_regfile_intregs_8__21_) );
  DFF_X2 decode_regfile_intregs_reg_8__22_ ( .D(n6460), .CK(clock), .Q(
        decode_regfile_intregs_8__22_) );
  DFF_X2 decode_regfile_intregs_reg_8__23_ ( .D(n6459), .CK(clock), .Q(
        decode_regfile_intregs_8__23_) );
  DFF_X2 decode_regfile_intregs_reg_8__24_ ( .D(n6458), .CK(clock), .Q(
        decode_regfile_intregs_8__24_) );
  DFF_X2 decode_regfile_intregs_reg_8__25_ ( .D(n6457), .CK(clock), .Q(
        decode_regfile_intregs_8__25_) );
  DFF_X2 decode_regfile_intregs_reg_8__26_ ( .D(n6456), .CK(clock), .Q(
        decode_regfile_intregs_8__26_) );
  DFF_X2 decode_regfile_intregs_reg_8__27_ ( .D(n6455), .CK(clock), .Q(
        decode_regfile_intregs_8__27_) );
  DFF_X2 decode_regfile_intregs_reg_8__28_ ( .D(n6454), .CK(clock), .Q(
        decode_regfile_intregs_8__28_) );
  DFF_X2 decode_regfile_intregs_reg_8__29_ ( .D(n6453), .CK(clock), .Q(
        decode_regfile_intregs_8__29_) );
  DFF_X2 decode_regfile_intregs_reg_8__30_ ( .D(n6452), .CK(clock), .Q(
        decode_regfile_intregs_8__30_) );
  DFF_X2 decode_regfile_intregs_reg_8__31_ ( .D(n6451), .CK(clock), .Q(
        decode_regfile_intregs_8__31_) );
  DFF_X2 decode_regfile_intregs_reg_7__0_ ( .D(n6450), .CK(clock), .Q(
        decode_regfile_intregs_7__0_) );
  DFF_X2 decode_regfile_intregs_reg_7__1_ ( .D(n6449), .CK(clock), .Q(
        decode_regfile_intregs_7__1_) );
  DFF_X2 decode_regfile_intregs_reg_7__2_ ( .D(n6448), .CK(clock), .Q(
        decode_regfile_intregs_7__2_) );
  DFF_X2 decode_regfile_intregs_reg_7__3_ ( .D(n6447), .CK(clock), .Q(
        decode_regfile_intregs_7__3_) );
  DFF_X2 decode_regfile_intregs_reg_7__4_ ( .D(n6446), .CK(clock), .Q(
        decode_regfile_intregs_7__4_) );
  DFF_X2 decode_regfile_intregs_reg_7__5_ ( .D(n6445), .CK(clock), .Q(
        decode_regfile_intregs_7__5_) );
  DFF_X2 decode_regfile_intregs_reg_7__6_ ( .D(n6444), .CK(clock), .Q(
        decode_regfile_intregs_7__6_) );
  DFF_X2 decode_regfile_intregs_reg_7__7_ ( .D(n6443), .CK(clock), .Q(
        decode_regfile_intregs_7__7_) );
  DFF_X2 decode_regfile_intregs_reg_7__8_ ( .D(n6442), .CK(clock), .Q(
        decode_regfile_intregs_7__8_) );
  DFF_X2 decode_regfile_intregs_reg_7__9_ ( .D(n6441), .CK(clock), .Q(
        decode_regfile_intregs_7__9_) );
  DFF_X2 decode_regfile_intregs_reg_7__10_ ( .D(n6440), .CK(clock), .Q(
        decode_regfile_intregs_7__10_) );
  DFF_X2 decode_regfile_intregs_reg_7__11_ ( .D(n6439), .CK(clock), .Q(
        decode_regfile_intregs_7__11_) );
  DFF_X2 decode_regfile_intregs_reg_7__12_ ( .D(n6438), .CK(clock), .Q(
        decode_regfile_intregs_7__12_) );
  DFF_X2 decode_regfile_intregs_reg_7__13_ ( .D(n6437), .CK(clock), .Q(
        decode_regfile_intregs_7__13_) );
  DFF_X2 decode_regfile_intregs_reg_7__14_ ( .D(n6436), .CK(clock), .Q(
        decode_regfile_intregs_7__14_) );
  DFF_X2 decode_regfile_intregs_reg_7__15_ ( .D(n6435), .CK(clock), .Q(
        decode_regfile_intregs_7__15_) );
  DFF_X2 decode_regfile_intregs_reg_7__16_ ( .D(n6434), .CK(clock), .Q(
        decode_regfile_intregs_7__16_) );
  DFF_X2 decode_regfile_intregs_reg_7__17_ ( .D(n6433), .CK(clock), .Q(
        decode_regfile_intregs_7__17_) );
  DFF_X2 decode_regfile_intregs_reg_7__18_ ( .D(n6432), .CK(clock), .Q(
        decode_regfile_intregs_7__18_) );
  DFF_X2 decode_regfile_intregs_reg_7__19_ ( .D(n6431), .CK(clock), .Q(
        decode_regfile_intregs_7__19_) );
  DFF_X2 decode_regfile_intregs_reg_7__20_ ( .D(n6430), .CK(clock), .Q(
        decode_regfile_intregs_7__20_) );
  DFF_X2 decode_regfile_intregs_reg_7__21_ ( .D(n6429), .CK(clock), .Q(
        decode_regfile_intregs_7__21_) );
  DFF_X2 decode_regfile_intregs_reg_7__22_ ( .D(n6428), .CK(clock), .Q(
        decode_regfile_intregs_7__22_) );
  DFF_X2 decode_regfile_intregs_reg_7__23_ ( .D(n6427), .CK(clock), .Q(
        decode_regfile_intregs_7__23_) );
  DFF_X2 decode_regfile_intregs_reg_7__24_ ( .D(n6426), .CK(clock), .Q(
        decode_regfile_intregs_7__24_) );
  DFF_X2 decode_regfile_intregs_reg_7__25_ ( .D(n6425), .CK(clock), .Q(
        decode_regfile_intregs_7__25_) );
  DFF_X2 decode_regfile_intregs_reg_7__26_ ( .D(n6424), .CK(clock), .Q(
        decode_regfile_intregs_7__26_) );
  DFF_X2 decode_regfile_intregs_reg_7__27_ ( .D(n6423), .CK(clock), .Q(
        decode_regfile_intregs_7__27_) );
  DFF_X2 decode_regfile_intregs_reg_7__28_ ( .D(n6422), .CK(clock), .Q(
        decode_regfile_intregs_7__28_) );
  DFF_X2 decode_regfile_intregs_reg_7__29_ ( .D(n6421), .CK(clock), .Q(
        decode_regfile_intregs_7__29_) );
  DFF_X2 decode_regfile_intregs_reg_7__30_ ( .D(n6420), .CK(clock), .Q(
        decode_regfile_intregs_7__30_) );
  DFF_X2 decode_regfile_intregs_reg_7__31_ ( .D(n6419), .CK(clock), .Q(
        decode_regfile_intregs_7__31_) );
  DFF_X2 decode_regfile_intregs_reg_6__0_ ( .D(n6418), .CK(clock), .Q(
        decode_regfile_intregs_6__0_) );
  DFF_X2 decode_regfile_intregs_reg_6__1_ ( .D(n6417), .CK(clock), .Q(
        decode_regfile_intregs_6__1_) );
  DFF_X2 decode_regfile_intregs_reg_6__2_ ( .D(n6416), .CK(clock), .Q(
        decode_regfile_intregs_6__2_) );
  DFF_X2 decode_regfile_intregs_reg_6__3_ ( .D(n6415), .CK(clock), .Q(
        decode_regfile_intregs_6__3_) );
  DFF_X2 decode_regfile_intregs_reg_6__4_ ( .D(n6414), .CK(clock), .Q(
        decode_regfile_intregs_6__4_) );
  DFF_X2 decode_regfile_intregs_reg_6__5_ ( .D(n6413), .CK(clock), .Q(
        decode_regfile_intregs_6__5_) );
  DFF_X2 decode_regfile_intregs_reg_6__6_ ( .D(n6412), .CK(clock), .Q(
        decode_regfile_intregs_6__6_) );
  DFF_X2 decode_regfile_intregs_reg_6__7_ ( .D(n6411), .CK(clock), .Q(
        decode_regfile_intregs_6__7_) );
  DFF_X2 decode_regfile_intregs_reg_6__8_ ( .D(n6410), .CK(clock), .Q(
        decode_regfile_intregs_6__8_) );
  DFF_X2 decode_regfile_intregs_reg_6__9_ ( .D(n6409), .CK(clock), .Q(
        decode_regfile_intregs_6__9_) );
  DFF_X2 decode_regfile_intregs_reg_6__10_ ( .D(n6408), .CK(clock), .Q(
        decode_regfile_intregs_6__10_) );
  DFF_X2 decode_regfile_intregs_reg_6__11_ ( .D(n6407), .CK(clock), .Q(
        decode_regfile_intregs_6__11_) );
  DFF_X2 decode_regfile_intregs_reg_6__12_ ( .D(n6406), .CK(clock), .Q(
        decode_regfile_intregs_6__12_) );
  DFF_X2 decode_regfile_intregs_reg_6__13_ ( .D(n6405), .CK(clock), .Q(
        decode_regfile_intregs_6__13_) );
  DFF_X2 decode_regfile_intregs_reg_6__14_ ( .D(n6404), .CK(clock), .Q(
        decode_regfile_intregs_6__14_) );
  DFF_X2 decode_regfile_intregs_reg_6__15_ ( .D(n6403), .CK(clock), .Q(
        decode_regfile_intregs_6__15_) );
  DFF_X2 decode_regfile_intregs_reg_6__16_ ( .D(n6402), .CK(clock), .Q(
        decode_regfile_intregs_6__16_) );
  DFF_X2 decode_regfile_intregs_reg_6__17_ ( .D(n6401), .CK(clock), .Q(
        decode_regfile_intregs_6__17_) );
  DFF_X2 decode_regfile_intregs_reg_6__18_ ( .D(n6400), .CK(clock), .Q(
        decode_regfile_intregs_6__18_) );
  DFF_X2 decode_regfile_intregs_reg_6__19_ ( .D(n6399), .CK(clock), .Q(
        decode_regfile_intregs_6__19_) );
  DFF_X2 decode_regfile_intregs_reg_6__20_ ( .D(n6398), .CK(clock), .Q(
        decode_regfile_intregs_6__20_) );
  DFF_X2 decode_regfile_intregs_reg_6__21_ ( .D(n6397), .CK(clock), .Q(
        decode_regfile_intregs_6__21_) );
  DFF_X2 decode_regfile_intregs_reg_6__22_ ( .D(n6396), .CK(clock), .Q(
        decode_regfile_intregs_6__22_) );
  DFF_X2 decode_regfile_intregs_reg_6__23_ ( .D(n6395), .CK(clock), .Q(
        decode_regfile_intregs_6__23_) );
  DFF_X2 decode_regfile_intregs_reg_6__24_ ( .D(n6394), .CK(clock), .Q(
        decode_regfile_intregs_6__24_) );
  DFF_X2 decode_regfile_intregs_reg_6__25_ ( .D(n6393), .CK(clock), .Q(
        decode_regfile_intregs_6__25_) );
  DFF_X2 decode_regfile_intregs_reg_6__26_ ( .D(n6392), .CK(clock), .Q(
        decode_regfile_intregs_6__26_) );
  DFF_X2 decode_regfile_intregs_reg_6__27_ ( .D(n6391), .CK(clock), .Q(
        decode_regfile_intregs_6__27_) );
  DFF_X2 decode_regfile_intregs_reg_6__28_ ( .D(n6390), .CK(clock), .Q(
        decode_regfile_intregs_6__28_) );
  DFF_X2 decode_regfile_intregs_reg_6__29_ ( .D(n6389), .CK(clock), .Q(
        decode_regfile_intregs_6__29_) );
  DFF_X2 decode_regfile_intregs_reg_6__30_ ( .D(n6388), .CK(clock), .Q(
        decode_regfile_intregs_6__30_) );
  DFF_X2 decode_regfile_intregs_reg_6__31_ ( .D(n6387), .CK(clock), .Q(
        decode_regfile_intregs_6__31_) );
  DFF_X2 decode_regfile_intregs_reg_5__0_ ( .D(n6386), .CK(clock), .Q(
        decode_regfile_intregs_5__0_) );
  DFF_X2 decode_regfile_intregs_reg_5__1_ ( .D(n6385), .CK(clock), .Q(
        decode_regfile_intregs_5__1_) );
  DFF_X2 decode_regfile_intregs_reg_5__2_ ( .D(n6384), .CK(clock), .Q(
        decode_regfile_intregs_5__2_) );
  DFF_X2 decode_regfile_intregs_reg_5__3_ ( .D(n6383), .CK(clock), .Q(
        decode_regfile_intregs_5__3_) );
  DFF_X2 decode_regfile_intregs_reg_5__4_ ( .D(n6382), .CK(clock), .Q(
        decode_regfile_intregs_5__4_) );
  DFF_X2 decode_regfile_intregs_reg_5__5_ ( .D(n6381), .CK(clock), .Q(
        decode_regfile_intregs_5__5_) );
  DFF_X2 decode_regfile_intregs_reg_5__6_ ( .D(n6380), .CK(clock), .Q(
        decode_regfile_intregs_5__6_) );
  DFF_X2 decode_regfile_intregs_reg_5__7_ ( .D(n6379), .CK(clock), .Q(
        decode_regfile_intregs_5__7_) );
  DFF_X2 decode_regfile_intregs_reg_5__8_ ( .D(n6378), .CK(clock), .Q(
        decode_regfile_intregs_5__8_) );
  DFF_X2 decode_regfile_intregs_reg_5__9_ ( .D(n6377), .CK(clock), .Q(
        decode_regfile_intregs_5__9_) );
  DFF_X2 decode_regfile_intregs_reg_5__10_ ( .D(n6376), .CK(clock), .Q(
        decode_regfile_intregs_5__10_) );
  DFF_X2 decode_regfile_intregs_reg_5__11_ ( .D(n6375), .CK(clock), .Q(
        decode_regfile_intregs_5__11_) );
  DFF_X2 decode_regfile_intregs_reg_5__12_ ( .D(n6374), .CK(clock), .Q(
        decode_regfile_intregs_5__12_) );
  DFF_X2 decode_regfile_intregs_reg_5__13_ ( .D(n6373), .CK(clock), .Q(
        decode_regfile_intregs_5__13_) );
  DFF_X2 decode_regfile_intregs_reg_5__14_ ( .D(n6372), .CK(clock), .Q(
        decode_regfile_intregs_5__14_) );
  DFF_X2 decode_regfile_intregs_reg_5__15_ ( .D(n6371), .CK(clock), .Q(
        decode_regfile_intregs_5__15_) );
  DFF_X2 decode_regfile_intregs_reg_5__16_ ( .D(n6370), .CK(clock), .Q(
        decode_regfile_intregs_5__16_) );
  DFF_X2 decode_regfile_intregs_reg_5__17_ ( .D(n6369), .CK(clock), .Q(
        decode_regfile_intregs_5__17_) );
  DFF_X2 decode_regfile_intregs_reg_5__18_ ( .D(n6368), .CK(clock), .Q(
        decode_regfile_intregs_5__18_) );
  DFF_X2 decode_regfile_intregs_reg_5__19_ ( .D(n6367), .CK(clock), .Q(
        decode_regfile_intregs_5__19_) );
  DFF_X2 decode_regfile_intregs_reg_5__20_ ( .D(n6366), .CK(clock), .Q(
        decode_regfile_intregs_5__20_) );
  DFF_X2 decode_regfile_intregs_reg_5__21_ ( .D(n6365), .CK(clock), .Q(
        decode_regfile_intregs_5__21_) );
  DFF_X2 decode_regfile_intregs_reg_5__22_ ( .D(n6364), .CK(clock), .Q(
        decode_regfile_intregs_5__22_) );
  DFF_X2 decode_regfile_intregs_reg_5__23_ ( .D(n6363), .CK(clock), .Q(
        decode_regfile_intregs_5__23_) );
  DFF_X2 decode_regfile_intregs_reg_5__24_ ( .D(n6362), .CK(clock), .Q(
        decode_regfile_intregs_5__24_) );
  DFF_X2 decode_regfile_intregs_reg_5__25_ ( .D(n6361), .CK(clock), .Q(
        decode_regfile_intregs_5__25_) );
  DFF_X2 decode_regfile_intregs_reg_5__26_ ( .D(n6360), .CK(clock), .Q(
        decode_regfile_intregs_5__26_) );
  DFF_X2 decode_regfile_intregs_reg_5__27_ ( .D(n6359), .CK(clock), .Q(
        decode_regfile_intregs_5__27_) );
  DFF_X2 decode_regfile_intregs_reg_5__28_ ( .D(n6358), .CK(clock), .Q(
        decode_regfile_intregs_5__28_) );
  DFF_X2 decode_regfile_intregs_reg_5__29_ ( .D(n6357), .CK(clock), .Q(
        decode_regfile_intregs_5__29_) );
  DFF_X2 decode_regfile_intregs_reg_5__30_ ( .D(n6356), .CK(clock), .Q(
        decode_regfile_intregs_5__30_) );
  DFF_X2 decode_regfile_intregs_reg_5__31_ ( .D(n6355), .CK(clock), .Q(
        decode_regfile_intregs_5__31_) );
  DFF_X2 decode_regfile_intregs_reg_4__0_ ( .D(n6354), .CK(clock), .Q(
        decode_regfile_intregs_4__0_) );
  DFF_X2 decode_regfile_intregs_reg_4__1_ ( .D(n6353), .CK(clock), .Q(
        decode_regfile_intregs_4__1_) );
  DFF_X2 decode_regfile_intregs_reg_4__2_ ( .D(n6352), .CK(clock), .Q(
        decode_regfile_intregs_4__2_) );
  DFF_X2 decode_regfile_intregs_reg_4__3_ ( .D(n6351), .CK(clock), .Q(
        decode_regfile_intregs_4__3_) );
  DFF_X2 decode_regfile_intregs_reg_4__4_ ( .D(n6350), .CK(clock), .Q(
        decode_regfile_intregs_4__4_) );
  DFF_X2 decode_regfile_intregs_reg_4__5_ ( .D(n6349), .CK(clock), .Q(
        decode_regfile_intregs_4__5_) );
  DFF_X2 decode_regfile_intregs_reg_4__6_ ( .D(n6348), .CK(clock), .Q(
        decode_regfile_intregs_4__6_) );
  DFF_X2 decode_regfile_intregs_reg_4__7_ ( .D(n6347), .CK(clock), .Q(
        decode_regfile_intregs_4__7_) );
  DFF_X2 decode_regfile_intregs_reg_4__8_ ( .D(n6346), .CK(clock), .Q(
        decode_regfile_intregs_4__8_) );
  DFF_X2 decode_regfile_intregs_reg_4__9_ ( .D(n6345), .CK(clock), .Q(
        decode_regfile_intregs_4__9_) );
  DFF_X2 decode_regfile_intregs_reg_4__10_ ( .D(n6344), .CK(clock), .Q(
        decode_regfile_intregs_4__10_) );
  DFF_X2 decode_regfile_intregs_reg_4__11_ ( .D(n6343), .CK(clock), .Q(
        decode_regfile_intregs_4__11_) );
  DFF_X2 decode_regfile_intregs_reg_4__12_ ( .D(n6342), .CK(clock), .Q(
        decode_regfile_intregs_4__12_) );
  DFF_X2 decode_regfile_intregs_reg_4__13_ ( .D(n6341), .CK(clock), .Q(
        decode_regfile_intregs_4__13_) );
  DFF_X2 decode_regfile_intregs_reg_4__14_ ( .D(n6340), .CK(clock), .Q(
        decode_regfile_intregs_4__14_) );
  DFF_X2 decode_regfile_intregs_reg_4__15_ ( .D(n6339), .CK(clock), .Q(
        decode_regfile_intregs_4__15_) );
  DFF_X2 decode_regfile_intregs_reg_4__16_ ( .D(n6338), .CK(clock), .Q(
        decode_regfile_intregs_4__16_) );
  DFF_X2 decode_regfile_intregs_reg_4__17_ ( .D(n6337), .CK(clock), .Q(
        decode_regfile_intregs_4__17_) );
  DFF_X2 decode_regfile_intregs_reg_4__18_ ( .D(n6336), .CK(clock), .Q(
        decode_regfile_intregs_4__18_) );
  DFF_X2 decode_regfile_intregs_reg_4__19_ ( .D(n6335), .CK(clock), .Q(
        decode_regfile_intregs_4__19_) );
  DFF_X2 decode_regfile_intregs_reg_4__20_ ( .D(n6334), .CK(clock), .Q(
        decode_regfile_intregs_4__20_) );
  DFF_X2 decode_regfile_intregs_reg_4__21_ ( .D(n6333), .CK(clock), .Q(
        decode_regfile_intregs_4__21_) );
  DFF_X2 decode_regfile_intregs_reg_4__22_ ( .D(n6332), .CK(clock), .Q(
        decode_regfile_intregs_4__22_) );
  DFF_X2 decode_regfile_intregs_reg_4__23_ ( .D(n6331), .CK(clock), .Q(
        decode_regfile_intregs_4__23_) );
  DFF_X2 decode_regfile_intregs_reg_4__24_ ( .D(n6330), .CK(clock), .Q(
        decode_regfile_intregs_4__24_) );
  DFF_X2 decode_regfile_intregs_reg_4__25_ ( .D(n6329), .CK(clock), .Q(
        decode_regfile_intregs_4__25_) );
  DFF_X2 decode_regfile_intregs_reg_4__26_ ( .D(n6328), .CK(clock), .Q(
        decode_regfile_intregs_4__26_) );
  DFF_X2 decode_regfile_intregs_reg_4__27_ ( .D(n6327), .CK(clock), .Q(
        decode_regfile_intregs_4__27_) );
  DFF_X2 decode_regfile_intregs_reg_4__28_ ( .D(n6326), .CK(clock), .Q(
        decode_regfile_intregs_4__28_) );
  DFF_X2 decode_regfile_intregs_reg_4__29_ ( .D(n6325), .CK(clock), .Q(
        decode_regfile_intregs_4__29_) );
  DFF_X2 decode_regfile_intregs_reg_4__30_ ( .D(n6324), .CK(clock), .Q(
        decode_regfile_intregs_4__30_) );
  DFF_X2 decode_regfile_intregs_reg_4__31_ ( .D(n6323), .CK(clock), .Q(
        decode_regfile_intregs_4__31_) );
  DFF_X2 decode_regfile_intregs_reg_3__0_ ( .D(n6322), .CK(clock), .Q(
        decode_regfile_intregs_3__0_) );
  DFF_X2 decode_regfile_intregs_reg_3__1_ ( .D(n6321), .CK(clock), .Q(
        decode_regfile_intregs_3__1_) );
  DFF_X2 decode_regfile_intregs_reg_3__2_ ( .D(n6320), .CK(clock), .Q(
        decode_regfile_intregs_3__2_) );
  DFF_X2 decode_regfile_intregs_reg_3__3_ ( .D(n6319), .CK(clock), .Q(
        decode_regfile_intregs_3__3_) );
  DFF_X2 decode_regfile_intregs_reg_3__4_ ( .D(n6318), .CK(clock), .Q(
        decode_regfile_intregs_3__4_) );
  DFF_X2 decode_regfile_intregs_reg_3__5_ ( .D(n6317), .CK(clock), .Q(
        decode_regfile_intregs_3__5_) );
  DFF_X2 decode_regfile_intregs_reg_3__6_ ( .D(n6316), .CK(clock), .Q(
        decode_regfile_intregs_3__6_) );
  DFF_X2 decode_regfile_intregs_reg_3__7_ ( .D(n6315), .CK(clock), .Q(
        decode_regfile_intregs_3__7_) );
  DFF_X2 decode_regfile_intregs_reg_3__8_ ( .D(n6314), .CK(clock), .Q(
        decode_regfile_intregs_3__8_) );
  DFF_X2 decode_regfile_intregs_reg_3__9_ ( .D(n6313), .CK(clock), .Q(
        decode_regfile_intregs_3__9_) );
  DFF_X2 decode_regfile_intregs_reg_3__10_ ( .D(n6312), .CK(clock), .Q(
        decode_regfile_intregs_3__10_) );
  DFF_X2 decode_regfile_intregs_reg_3__11_ ( .D(n6311), .CK(clock), .Q(
        decode_regfile_intregs_3__11_) );
  DFF_X2 decode_regfile_intregs_reg_3__12_ ( .D(n6310), .CK(clock), .Q(
        decode_regfile_intregs_3__12_) );
  DFF_X2 decode_regfile_intregs_reg_3__13_ ( .D(n6309), .CK(clock), .Q(
        decode_regfile_intregs_3__13_) );
  DFF_X2 decode_regfile_intregs_reg_3__14_ ( .D(n6308), .CK(clock), .Q(
        decode_regfile_intregs_3__14_) );
  DFF_X2 decode_regfile_intregs_reg_3__15_ ( .D(n6307), .CK(clock), .Q(
        decode_regfile_intregs_3__15_) );
  DFF_X2 decode_regfile_intregs_reg_3__16_ ( .D(n6306), .CK(clock), .Q(
        decode_regfile_intregs_3__16_) );
  DFF_X2 decode_regfile_intregs_reg_3__17_ ( .D(n6305), .CK(clock), .Q(
        decode_regfile_intregs_3__17_) );
  DFF_X2 decode_regfile_intregs_reg_3__18_ ( .D(n6304), .CK(clock), .Q(
        decode_regfile_intregs_3__18_) );
  DFF_X2 decode_regfile_intregs_reg_3__19_ ( .D(n6303), .CK(clock), .Q(
        decode_regfile_intregs_3__19_) );
  DFF_X2 decode_regfile_intregs_reg_3__20_ ( .D(n6302), .CK(clock), .Q(
        decode_regfile_intregs_3__20_) );
  DFF_X2 decode_regfile_intregs_reg_3__21_ ( .D(n6301), .CK(clock), .Q(
        decode_regfile_intregs_3__21_) );
  DFF_X2 decode_regfile_intregs_reg_3__22_ ( .D(n6300), .CK(clock), .Q(
        decode_regfile_intregs_3__22_) );
  DFF_X2 decode_regfile_intregs_reg_3__23_ ( .D(n6299), .CK(clock), .Q(
        decode_regfile_intregs_3__23_) );
  DFF_X2 decode_regfile_intregs_reg_3__24_ ( .D(n6298), .CK(clock), .Q(
        decode_regfile_intregs_3__24_) );
  DFF_X2 decode_regfile_intregs_reg_3__25_ ( .D(n6297), .CK(clock), .Q(
        decode_regfile_intregs_3__25_) );
  DFF_X2 decode_regfile_intregs_reg_3__26_ ( .D(n6296), .CK(clock), .Q(
        decode_regfile_intregs_3__26_) );
  DFF_X2 decode_regfile_intregs_reg_3__27_ ( .D(n6295), .CK(clock), .Q(
        decode_regfile_intregs_3__27_) );
  DFF_X2 decode_regfile_intregs_reg_3__28_ ( .D(n6294), .CK(clock), .Q(
        decode_regfile_intregs_3__28_) );
  DFF_X2 decode_regfile_intregs_reg_3__29_ ( .D(n6293), .CK(clock), .Q(
        decode_regfile_intregs_3__29_) );
  DFF_X2 decode_regfile_intregs_reg_3__30_ ( .D(n6292), .CK(clock), .Q(
        decode_regfile_intregs_3__30_) );
  DFF_X2 decode_regfile_intregs_reg_3__31_ ( .D(n6291), .CK(clock), .Q(
        decode_regfile_intregs_3__31_) );
  DFF_X2 decode_regfile_intregs_reg_2__0_ ( .D(n6290), .CK(clock), .Q(
        decode_regfile_intregs_2__0_) );
  DFF_X2 decode_regfile_intregs_reg_2__1_ ( .D(n6289), .CK(clock), .Q(
        decode_regfile_intregs_2__1_) );
  DFF_X2 decode_regfile_intregs_reg_2__2_ ( .D(n6288), .CK(clock), .Q(
        decode_regfile_intregs_2__2_) );
  DFF_X2 decode_regfile_intregs_reg_2__3_ ( .D(n6287), .CK(clock), .Q(
        decode_regfile_intregs_2__3_) );
  DFF_X2 decode_regfile_intregs_reg_2__4_ ( .D(n6286), .CK(clock), .Q(
        decode_regfile_intregs_2__4_) );
  DFF_X2 decode_regfile_intregs_reg_2__5_ ( .D(n6285), .CK(clock), .Q(
        decode_regfile_intregs_2__5_) );
  DFF_X2 decode_regfile_intregs_reg_2__6_ ( .D(n6284), .CK(clock), .Q(
        decode_regfile_intregs_2__6_) );
  DFF_X2 decode_regfile_intregs_reg_2__7_ ( .D(n6283), .CK(clock), .Q(
        decode_regfile_intregs_2__7_) );
  DFF_X2 decode_regfile_intregs_reg_2__8_ ( .D(n6282), .CK(clock), .Q(
        decode_regfile_intregs_2__8_) );
  DFF_X2 decode_regfile_intregs_reg_2__9_ ( .D(n6281), .CK(clock), .Q(
        decode_regfile_intregs_2__9_) );
  DFF_X2 decode_regfile_intregs_reg_2__10_ ( .D(n6280), .CK(clock), .Q(
        decode_regfile_intregs_2__10_) );
  DFF_X2 decode_regfile_intregs_reg_2__11_ ( .D(n6279), .CK(clock), .Q(
        decode_regfile_intregs_2__11_) );
  DFF_X2 decode_regfile_intregs_reg_2__12_ ( .D(n6278), .CK(clock), .Q(
        decode_regfile_intregs_2__12_) );
  DFF_X2 decode_regfile_intregs_reg_2__13_ ( .D(n6277), .CK(clock), .Q(
        decode_regfile_intregs_2__13_) );
  DFF_X2 decode_regfile_intregs_reg_2__14_ ( .D(n6276), .CK(clock), .Q(
        decode_regfile_intregs_2__14_) );
  DFF_X2 decode_regfile_intregs_reg_2__15_ ( .D(n6275), .CK(clock), .Q(
        decode_regfile_intregs_2__15_) );
  DFF_X2 decode_regfile_intregs_reg_2__16_ ( .D(n6274), .CK(clock), .Q(
        decode_regfile_intregs_2__16_) );
  DFF_X2 decode_regfile_intregs_reg_2__17_ ( .D(n6273), .CK(clock), .Q(
        decode_regfile_intregs_2__17_) );
  DFF_X2 decode_regfile_intregs_reg_2__18_ ( .D(n6272), .CK(clock), .Q(
        decode_regfile_intregs_2__18_) );
  DFF_X2 decode_regfile_intregs_reg_2__19_ ( .D(n6271), .CK(clock), .Q(
        decode_regfile_intregs_2__19_) );
  DFF_X2 decode_regfile_intregs_reg_2__20_ ( .D(n6270), .CK(clock), .Q(
        decode_regfile_intregs_2__20_) );
  DFF_X2 decode_regfile_intregs_reg_2__21_ ( .D(n6269), .CK(clock), .Q(
        decode_regfile_intregs_2__21_) );
  DFF_X2 decode_regfile_intregs_reg_2__22_ ( .D(n6268), .CK(clock), .Q(
        decode_regfile_intregs_2__22_) );
  DFF_X2 decode_regfile_intregs_reg_2__23_ ( .D(n6267), .CK(clock), .Q(
        decode_regfile_intregs_2__23_) );
  DFF_X2 decode_regfile_intregs_reg_2__24_ ( .D(n6266), .CK(clock), .Q(
        decode_regfile_intregs_2__24_) );
  DFF_X2 decode_regfile_intregs_reg_2__25_ ( .D(n6265), .CK(clock), .Q(
        decode_regfile_intregs_2__25_) );
  DFF_X2 decode_regfile_intregs_reg_2__26_ ( .D(n6264), .CK(clock), .Q(
        decode_regfile_intregs_2__26_) );
  DFF_X2 decode_regfile_intregs_reg_2__27_ ( .D(n6263), .CK(clock), .Q(
        decode_regfile_intregs_2__27_) );
  DFF_X2 decode_regfile_intregs_reg_2__28_ ( .D(n6262), .CK(clock), .Q(
        decode_regfile_intregs_2__28_) );
  DFF_X2 decode_regfile_intregs_reg_2__29_ ( .D(n6261), .CK(clock), .Q(
        decode_regfile_intregs_2__29_) );
  DFF_X2 decode_regfile_intregs_reg_2__30_ ( .D(n6260), .CK(clock), .Q(
        decode_regfile_intregs_2__30_) );
  DFF_X2 decode_regfile_intregs_reg_2__31_ ( .D(n6259), .CK(clock), .Q(
        decode_regfile_intregs_2__31_) );
  DFF_X2 decode_regfile_intregs_reg_1__0_ ( .D(n6258), .CK(clock), .Q(
        decode_regfile_intregs_1__0_) );
  DFF_X2 decode_regfile_intregs_reg_1__1_ ( .D(n6257), .CK(clock), .Q(
        decode_regfile_intregs_1__1_) );
  DFF_X2 decode_regfile_intregs_reg_1__2_ ( .D(n6256), .CK(clock), .Q(
        decode_regfile_intregs_1__2_) );
  DFF_X2 decode_regfile_intregs_reg_1__3_ ( .D(n6255), .CK(clock), .Q(
        decode_regfile_intregs_1__3_) );
  DFF_X2 decode_regfile_intregs_reg_1__4_ ( .D(n6254), .CK(clock), .Q(
        decode_regfile_intregs_1__4_) );
  DFF_X2 decode_regfile_intregs_reg_1__5_ ( .D(n6253), .CK(clock), .Q(
        decode_regfile_intregs_1__5_) );
  DFF_X2 decode_regfile_intregs_reg_1__6_ ( .D(n6252), .CK(clock), .Q(
        decode_regfile_intregs_1__6_) );
  DFF_X2 decode_regfile_intregs_reg_1__7_ ( .D(n6251), .CK(clock), .Q(
        decode_regfile_intregs_1__7_) );
  DFF_X2 decode_regfile_intregs_reg_1__8_ ( .D(n6250), .CK(clock), .Q(
        decode_regfile_intregs_1__8_) );
  DFF_X2 decode_regfile_intregs_reg_1__9_ ( .D(n6249), .CK(clock), .Q(
        decode_regfile_intregs_1__9_) );
  DFF_X2 decode_regfile_intregs_reg_1__10_ ( .D(n6248), .CK(clock), .Q(
        decode_regfile_intregs_1__10_) );
  DFF_X2 decode_regfile_intregs_reg_1__11_ ( .D(n6247), .CK(clock), .Q(
        decode_regfile_intregs_1__11_) );
  DFF_X2 decode_regfile_intregs_reg_1__12_ ( .D(n6246), .CK(clock), .Q(
        decode_regfile_intregs_1__12_) );
  DFF_X2 decode_regfile_intregs_reg_1__13_ ( .D(n6245), .CK(clock), .Q(
        decode_regfile_intregs_1__13_) );
  DFF_X2 decode_regfile_intregs_reg_1__14_ ( .D(n6244), .CK(clock), .Q(
        decode_regfile_intregs_1__14_) );
  DFF_X2 decode_regfile_intregs_reg_1__15_ ( .D(n6243), .CK(clock), .Q(
        decode_regfile_intregs_1__15_) );
  DFF_X2 decode_regfile_intregs_reg_1__16_ ( .D(n6242), .CK(clock), .Q(
        decode_regfile_intregs_1__16_) );
  DFF_X2 decode_regfile_intregs_reg_1__17_ ( .D(n6241), .CK(clock), .Q(
        decode_regfile_intregs_1__17_) );
  DFF_X2 decode_regfile_intregs_reg_1__18_ ( .D(n6240), .CK(clock), .Q(
        decode_regfile_intregs_1__18_) );
  DFF_X2 decode_regfile_intregs_reg_1__19_ ( .D(n6239), .CK(clock), .Q(
        decode_regfile_intregs_1__19_) );
  DFF_X2 decode_regfile_intregs_reg_1__20_ ( .D(n6238), .CK(clock), .Q(
        decode_regfile_intregs_1__20_) );
  DFF_X2 decode_regfile_intregs_reg_1__21_ ( .D(n6237), .CK(clock), .Q(
        decode_regfile_intregs_1__21_) );
  DFF_X2 decode_regfile_intregs_reg_1__22_ ( .D(n6236), .CK(clock), .Q(
        decode_regfile_intregs_1__22_) );
  DFF_X2 decode_regfile_intregs_reg_1__23_ ( .D(n6235), .CK(clock), .Q(
        decode_regfile_intregs_1__23_) );
  DFF_X2 decode_regfile_intregs_reg_1__24_ ( .D(n6234), .CK(clock), .Q(
        decode_regfile_intregs_1__24_) );
  DFF_X2 decode_regfile_intregs_reg_1__25_ ( .D(n6233), .CK(clock), .Q(
        decode_regfile_intregs_1__25_) );
  DFF_X2 decode_regfile_intregs_reg_1__26_ ( .D(n6232), .CK(clock), .Q(
        decode_regfile_intregs_1__26_) );
  DFF_X2 decode_regfile_intregs_reg_1__27_ ( .D(n6231), .CK(clock), .Q(
        decode_regfile_intregs_1__27_) );
  DFF_X2 decode_regfile_intregs_reg_1__28_ ( .D(n6230), .CK(clock), .Q(
        decode_regfile_intregs_1__28_) );
  DFF_X2 decode_regfile_intregs_reg_1__29_ ( .D(n6229), .CK(clock), .Q(
        decode_regfile_intregs_1__29_) );
  DFF_X2 decode_regfile_intregs_reg_1__30_ ( .D(n6228), .CK(clock), .Q(
        decode_regfile_intregs_1__30_) );
  DFF_X2 decode_regfile_intregs_reg_1__31_ ( .D(n6227), .CK(clock), .Q(
        decode_regfile_intregs_1__31_) );
  DFF_X2 decode_regfile_intregs_reg_0__0_ ( .D(n6226), .CK(clock), .Q(
        decode_regfile_intregs_0__0_) );
  DFF_X2 decode_regfile_intregs_reg_0__1_ ( .D(n6225), .CK(clock), .Q(
        decode_regfile_intregs_0__1_) );
  DFF_X2 decode_regfile_intregs_reg_0__2_ ( .D(n6224), .CK(clock), .Q(
        decode_regfile_intregs_0__2_) );
  DFF_X2 decode_regfile_intregs_reg_0__3_ ( .D(n6223), .CK(clock), .Q(
        decode_regfile_intregs_0__3_) );
  DFF_X2 decode_regfile_intregs_reg_0__4_ ( .D(n6222), .CK(clock), .Q(
        decode_regfile_intregs_0__4_) );
  DFF_X2 decode_regfile_intregs_reg_0__5_ ( .D(n6221), .CK(clock), .Q(
        decode_regfile_intregs_0__5_) );
  DFF_X2 decode_regfile_intregs_reg_0__6_ ( .D(n6220), .CK(clock), .Q(
        decode_regfile_intregs_0__6_) );
  DFF_X2 decode_regfile_intregs_reg_0__7_ ( .D(n6219), .CK(clock), .Q(
        decode_regfile_intregs_0__7_) );
  DFF_X2 decode_regfile_intregs_reg_0__8_ ( .D(n6218), .CK(clock), .Q(
        decode_regfile_intregs_0__8_) );
  DFF_X2 decode_regfile_intregs_reg_0__9_ ( .D(n6217), .CK(clock), .Q(
        decode_regfile_intregs_0__9_) );
  DFF_X2 decode_regfile_intregs_reg_0__10_ ( .D(n6216), .CK(clock), .Q(
        decode_regfile_intregs_0__10_) );
  DFF_X2 decode_regfile_intregs_reg_0__11_ ( .D(n6215), .CK(clock), .Q(
        decode_regfile_intregs_0__11_) );
  DFF_X2 decode_regfile_intregs_reg_0__12_ ( .D(n6214), .CK(clock), .Q(
        decode_regfile_intregs_0__12_) );
  DFF_X2 decode_regfile_intregs_reg_0__13_ ( .D(n6213), .CK(clock), .Q(
        decode_regfile_intregs_0__13_) );
  DFF_X2 decode_regfile_intregs_reg_0__14_ ( .D(n6212), .CK(clock), .Q(
        decode_regfile_intregs_0__14_) );
  DFF_X2 decode_regfile_intregs_reg_0__15_ ( .D(n6211), .CK(clock), .Q(
        decode_regfile_intregs_0__15_) );
  DFF_X2 decode_regfile_intregs_reg_0__16_ ( .D(n6210), .CK(clock), .Q(
        decode_regfile_intregs_0__16_) );
  DFF_X2 decode_regfile_intregs_reg_0__17_ ( .D(n6209), .CK(clock), .Q(
        decode_regfile_intregs_0__17_) );
  DFF_X2 decode_regfile_intregs_reg_0__18_ ( .D(n6208), .CK(clock), .Q(
        decode_regfile_intregs_0__18_) );
  DFF_X2 decode_regfile_intregs_reg_0__19_ ( .D(n6207), .CK(clock), .Q(
        decode_regfile_intregs_0__19_) );
  DFF_X2 decode_regfile_intregs_reg_0__20_ ( .D(n6206), .CK(clock), .Q(
        decode_regfile_intregs_0__20_) );
  DFF_X2 decode_regfile_intregs_reg_0__21_ ( .D(n6205), .CK(clock), .Q(
        decode_regfile_intregs_0__21_) );
  DFF_X2 decode_regfile_intregs_reg_0__22_ ( .D(n6204), .CK(clock), .Q(
        decode_regfile_intregs_0__22_) );
  DFF_X2 decode_regfile_intregs_reg_0__23_ ( .D(n6203), .CK(clock), .Q(
        decode_regfile_intregs_0__23_) );
  DFF_X2 decode_regfile_intregs_reg_0__24_ ( .D(n6202), .CK(clock), .Q(
        decode_regfile_intregs_0__24_) );
  DFF_X2 decode_regfile_intregs_reg_0__25_ ( .D(n6201), .CK(clock), .Q(
        decode_regfile_intregs_0__25_) );
  DFF_X2 decode_regfile_intregs_reg_0__26_ ( .D(n6200), .CK(clock), .Q(
        decode_regfile_intregs_0__26_) );
  DFF_X2 decode_regfile_intregs_reg_0__27_ ( .D(n6199), .CK(clock), .Q(
        decode_regfile_intregs_0__27_) );
  DFF_X2 decode_regfile_intregs_reg_0__28_ ( .D(n6198), .CK(clock), .Q(
        decode_regfile_intregs_0__28_) );
  DFF_X2 decode_regfile_intregs_reg_0__29_ ( .D(n6197), .CK(clock), .Q(
        decode_regfile_intregs_0__29_) );
  DFF_X2 decode_regfile_intregs_reg_0__30_ ( .D(n6196), .CK(clock), .Q(
        decode_regfile_intregs_0__30_) );
  DFF_X2 decode_regfile_intregs_reg_0__31_ ( .D(n6195), .CK(clock), .Q(
        decode_regfile_intregs_0__31_) );
  OAI221_X2 U48 ( .B1(n13776), .B2(n38), .C1(n16296), .C2(n13775), .A(n57), 
        .ZN(execstage_register_N99) );
  OAI221_X2 U50 ( .B1(n13776), .B2(n37), .C1(n16294), .C2(n13775), .A(n63), 
        .ZN(execstage_register_N98) );
  OAI221_X2 U52 ( .B1(n13776), .B2(n36), .C1(n16312), .C2(n13775), .A(n66), 
        .ZN(execstage_register_N97) );
  OAI221_X2 U54 ( .B1(n13776), .B2(n35), .C1(n16313), .C2(n13775), .A(n69), 
        .ZN(execstage_register_N96) );
  OAI221_X2 U56 ( .B1(n13776), .B2(n34), .C1(n16311), .C2(n13775), .A(n72), 
        .ZN(execstage_register_N95) );
  OAI221_X2 U58 ( .B1(n13776), .B2(n33), .C1(n16316), .C2(n13775), .A(n75), 
        .ZN(execstage_register_N94) );
  OAI221_X2 U60 ( .B1(n13776), .B2(n32), .C1(n16319), .C2(n13775), .A(n78), 
        .ZN(execstage_register_N93) );
  OAI221_X2 U62 ( .B1(n13776), .B2(n31), .C1(n16256), .C2(n13775), .A(n81), 
        .ZN(execstage_register_N92) );
  OAI221_X2 U64 ( .B1(n13776), .B2(n30), .C1(n16324), .C2(n13775), .A(n84), 
        .ZN(execstage_register_N91) );
  OAI221_X2 U66 ( .B1(n13776), .B2(n29), .C1(n16349), .C2(n13775), .A(n87), 
        .ZN(execstage_register_N90) );
  AND2_X2 U68 ( .A1(aluctrl_0[0]), .A2(n13809), .ZN(execstage_register_N9) );
  OAI221_X2 U69 ( .B1(n13776), .B2(n28), .C1(n16352), .C2(n13774), .A(n91), 
        .ZN(execstage_register_N89) );
  OAI221_X2 U71 ( .B1(n13777), .B2(n27), .C1(n16333), .C2(n13774), .A(n94), 
        .ZN(execstage_register_N88) );
  OAI221_X2 U73 ( .B1(n13777), .B2(n26), .C1(n16403), .C2(n13774), .A(n97), 
        .ZN(execstage_register_N87) );
  OAI221_X2 U75 ( .B1(n13777), .B2(n25), .C1(n16387), .C2(n13774), .A(n100), 
        .ZN(execstage_register_N86) );
  OAI221_X2 U77 ( .B1(n13777), .B2(n24), .C1(n16400), .C2(n13774), .A(n103), 
        .ZN(execstage_register_N85) );
  OAI221_X2 U79 ( .B1(n13777), .B2(n23), .C1(n16397), .C2(n13774), .A(n106), 
        .ZN(execstage_register_N84) );
  OAI221_X2 U81 ( .B1(n13777), .B2(n22), .C1(n16212), .C2(n13774), .A(n109), 
        .ZN(execstage_register_N83) );
  AND2_X2 U83 ( .A1(n13809), .A2(n111), .ZN(execstage_register_N82) );
  AND2_X2 U84 ( .A1(n13809), .A2(n112), .ZN(execstage_register_N81) );
  AND2_X2 U85 ( .A1(n13809), .A2(n113), .ZN(execstage_register_N80) );
  AND2_X2 U86 ( .A1(n13803), .A2(n114), .ZN(execstage_register_N79) );
  AND2_X2 U87 ( .A1(n13809), .A2(n115), .ZN(execstage_register_N78) );
  AND2_X2 U88 ( .A1(n13809), .A2(n116), .ZN(execstage_register_N77) );
  AND2_X2 U89 ( .A1(n13809), .A2(n117), .ZN(execstage_register_N76) );
  AND2_X2 U90 ( .A1(n13809), .A2(n118), .ZN(execstage_register_N75) );
  AND2_X2 U91 ( .A1(n13809), .A2(n119), .ZN(execstage_register_N74) );
  AND2_X2 U92 ( .A1(n13809), .A2(n120), .ZN(execstage_register_N73) );
  OR4_X2 U110 ( .A1(n8749), .A2(n147), .A3(n148), .A4(imm32_0[5]), .ZN(n139)
         );
  AND2_X2 U138 ( .A1(jal_0), .A2(n13809), .ZN(execstage_register_N18) );
  NOR4_X2 U153 ( .A1(imm32_0[1]), .A2(n8748), .A3(n191), .A4(n20), .ZN(
        execstage_register_N14) );
  NAND2_X2 U165 ( .A1(imm32_0[5]), .A2(n13809), .ZN(n20) );
  OR3_X2 U166 ( .A1(n8749), .A2(n147), .A3(n16588), .ZN(n191) );
  AND2_X2 U177 ( .A1(aluctrl_0[3]), .A2(n13809), .ZN(execstage_register_N12)
         );
  OAI221_X2 U178 ( .B1(n10955), .B2(n215), .C1(n149), .C2(n19), .A(n135), .ZN(
        execstage_register_N119) );
  NAND2_X2 U179 ( .A1(imm32_0[15]), .A2(n13809), .ZN(n19) );
  OAI221_X2 U181 ( .B1(n10943), .B2(n215), .C1(n149), .C2(n18), .A(n135), .ZN(
        execstage_register_N118) );
  NAND2_X2 U182 ( .A1(imm32_0[14]), .A2(n13809), .ZN(n18) );
  OAI221_X2 U184 ( .B1(n13799), .B2(n215), .C1(n149), .C2(n17), .A(n135), .ZN(
        execstage_register_N117) );
  NAND2_X2 U185 ( .A1(imm32_0[13]), .A2(n13809), .ZN(n17) );
  OAI221_X2 U187 ( .B1(n13800), .B2(n215), .C1(n149), .C2(n16), .A(n135), .ZN(
        execstage_register_N116) );
  NAND2_X2 U188 ( .A1(imm32_0[12]), .A2(n13809), .ZN(n16) );
  OAI221_X2 U190 ( .B1(n13802), .B2(n215), .C1(n149), .C2(n15), .A(n135), .ZN(
        execstage_register_N115) );
  OR2_X2 U191 ( .A1(n220), .A2(n13808), .ZN(n135) );
  NAND2_X2 U192 ( .A1(imm32_0[11]), .A2(n13809), .ZN(n15) );
  NAND2_X2 U193 ( .A1(n13809), .A2(n149), .ZN(n215) );
  OAI221_X2 U195 ( .B1(n13777), .B2(n53), .C1(n16176), .C2(n13774), .A(n222), 
        .ZN(execstage_register_N114) );
  OAI221_X2 U197 ( .B1(n13777), .B2(n52), .C1(n16177), .C2(n13774), .A(n225), 
        .ZN(execstage_register_N113) );
  OAI221_X2 U199 ( .B1(n13777), .B2(n51), .C1(n16180), .C2(n13774), .A(n228), 
        .ZN(execstage_register_N112) );
  OAI221_X2 U201 ( .B1(n13777), .B2(n50), .C1(n16179), .C2(n13774), .A(n231), 
        .ZN(execstage_register_N111) );
  OAI221_X2 U203 ( .B1(n13777), .B2(n49), .C1(n16178), .C2(n13773), .A(n234), 
        .ZN(execstage_register_N110) );
  AND2_X2 U205 ( .A1(aluctrl_0[2]), .A2(n13809), .ZN(execstage_register_N11)
         );
  OAI221_X2 U206 ( .B1(n13778), .B2(n48), .C1(n16190), .C2(n13773), .A(n237), 
        .ZN(execstage_register_N109) );
  OAI221_X2 U208 ( .B1(n13778), .B2(n47), .C1(n16189), .C2(n13773), .A(n240), 
        .ZN(execstage_register_N108) );
  OAI221_X2 U210 ( .B1(n13778), .B2(n46), .C1(n16197), .C2(n13773), .A(n243), 
        .ZN(execstage_register_N107) );
  OAI221_X2 U212 ( .B1(n13778), .B2(n45), .C1(n16196), .C2(n13773), .A(n246), 
        .ZN(execstage_register_N106) );
  OAI221_X2 U214 ( .B1(n13778), .B2(n44), .C1(n16195), .C2(n13773), .A(n249), 
        .ZN(execstage_register_N105) );
  OAI221_X2 U216 ( .B1(n13778), .B2(n43), .C1(n16194), .C2(n13773), .A(n252), 
        .ZN(execstage_register_N104) );
  OAI221_X2 U218 ( .B1(n13778), .B2(n42), .C1(n16193), .C2(n13773), .A(n255), 
        .ZN(execstage_register_N103) );
  OAI221_X2 U220 ( .B1(n13778), .B2(n41), .C1(n16209), .C2(n13773), .A(n258), 
        .ZN(execstage_register_N102) );
  OAI221_X2 U222 ( .B1(n13778), .B2(n40), .C1(n16210), .C2(n13773), .A(n261), 
        .ZN(execstage_register_N101) );
  OAI221_X2 U224 ( .B1(n13778), .B2(n39), .C1(n16211), .C2(n13773), .A(n264), 
        .ZN(execstage_register_N100) );
  AND2_X2 U234 ( .A1(aluctrl_0[1]), .A2(n13809), .ZN(execstage_register_N10)
         );
  AND4_X2 U240 ( .A1(n16591), .A2(n277), .A3(n278), .A4(n279), .ZN(n162) );
  AND4_X2 U241 ( .A1(n280), .A2(n281), .A3(n282), .A4(n283), .ZN(n279) );
  AND3_X2 U248 ( .A1(n142), .A2(n282), .A3(n159), .ZN(n286) );
  AND4_X2 U249 ( .A1(n161), .A2(n292), .A3(n293), .A4(n294), .ZN(n159) );
  NAND4_X2 U251 ( .A1(n16600), .A2(n16591), .A3(n299), .A4(n300), .ZN(n145) );
  AND4_X2 U252 ( .A1(n280), .A2(n281), .A3(n301), .A4(n302), .ZN(n300) );
  NAND2_X2 U373 ( .A1(n16592), .A2(n320), .ZN(n312) );
  XOR2_X2 U374 ( .A(n8716), .B(n321), .Z(n320) );
  NAND4_X2 U375 ( .A1(n322), .A2(n323), .A3(n324), .A4(n325), .ZN(n321) );
  NOR4_X2 U376 ( .A1(n326), .A2(n327), .A3(n328), .A4(n329), .ZN(n325) );
  NAND4_X2 U377 ( .A1(n16170), .A2(n16171), .A3(n16172), .A4(n16173), .ZN(n329) );
  OAI221_X2 U379 ( .B1(n16311), .B2(n13758), .C1(n34), .C2(n13755), .A(n333), 
        .ZN(n330) );
  NAND2_X2 U381 ( .A1(mem_ExecResult[12]), .A2(n8725), .ZN(n34) );
  OAI221_X2 U384 ( .B1(n16313), .B2(n13758), .C1(n35), .C2(n13756), .A(n339), 
        .ZN(n338) );
  NAND2_X2 U386 ( .A1(mem_ExecResult[13]), .A2(n8725), .ZN(n35) );
  OAI221_X2 U389 ( .B1(n16312), .B2(n13758), .C1(n36), .C2(n13756), .A(n341), 
        .ZN(n340) );
  NAND2_X2 U391 ( .A1(mem_ExecResult[14]), .A2(n8725), .ZN(n36) );
  OAI221_X2 U394 ( .B1(n16294), .B2(n13758), .C1(n37), .C2(n13756), .A(n343), 
        .ZN(n342) );
  NAND2_X2 U396 ( .A1(mem_ExecResult[15]), .A2(n8725), .ZN(n37) );
  NAND4_X2 U398 ( .A1(n16166), .A2(n16167), .A3(n16168), .A4(n16169), .ZN(n328) );
  OAI221_X2 U400 ( .B1(n16324), .B2(n13758), .C1(n30), .C2(n13756), .A(n345), 
        .ZN(n344) );
  NAND2_X2 U402 ( .A1(mem_ExecResult[8]), .A2(n8725), .ZN(n30) );
  OAI221_X2 U405 ( .B1(n16256), .B2(n13758), .C1(n31), .C2(n13756), .A(n347), 
        .ZN(n346) );
  NAND2_X2 U407 ( .A1(mem_ExecResult[9]), .A2(n8725), .ZN(n31) );
  OAI221_X2 U410 ( .B1(n16319), .B2(n13758), .C1(n32), .C2(n13756), .A(n349), 
        .ZN(n348) );
  NAND2_X2 U412 ( .A1(mem_ExecResult[10]), .A2(n8725), .ZN(n32) );
  OAI221_X2 U415 ( .B1(n16316), .B2(n13758), .C1(n33), .C2(n13755), .A(n351), 
        .ZN(n350) );
  NAND2_X2 U417 ( .A1(mem_ExecResult[11]), .A2(n8725), .ZN(n33) );
  NAND4_X2 U419 ( .A1(n16162), .A2(n16163), .A3(n16164), .A4(n16165), .ZN(n327) );
  OAI221_X2 U421 ( .B1(n16403), .B2(n13758), .C1(n26), .C2(n13755), .A(n353), 
        .ZN(n352) );
  NAND2_X2 U423 ( .A1(mem_ExecResult[4]), .A2(n8725), .ZN(n26) );
  OAI221_X2 U426 ( .B1(n16333), .B2(n13758), .C1(n27), .C2(n13755), .A(n355), 
        .ZN(n354) );
  NAND2_X2 U428 ( .A1(mem_ExecResult[5]), .A2(n8725), .ZN(n27) );
  OAI221_X2 U431 ( .B1(n16352), .B2(n13758), .C1(n28), .C2(n13755), .A(n357), 
        .ZN(n356) );
  NAND2_X2 U433 ( .A1(mem_ExecResult[6]), .A2(n13127), .ZN(n28) );
  OAI221_X2 U436 ( .B1(n16349), .B2(n13759), .C1(n29), .C2(n13755), .A(n359), 
        .ZN(n358) );
  NAND2_X2 U438 ( .A1(mem_ExecResult[7]), .A2(n13127), .ZN(n29) );
  NAND4_X2 U440 ( .A1(n16158), .A2(n16159), .A3(n16160), .A4(n16161), .ZN(n326) );
  OAI221_X2 U442 ( .B1(n16212), .B2(n13759), .C1(n22), .C2(n13755), .A(n361), 
        .ZN(n360) );
  NAND2_X2 U444 ( .A1(mem_ExecResult[0]), .A2(n13127), .ZN(n22) );
  OAI221_X2 U447 ( .B1(n16397), .B2(n13759), .C1(n23), .C2(n13755), .A(n363), 
        .ZN(n362) );
  NAND2_X2 U449 ( .A1(mem_ExecResult[1]), .A2(n13127), .ZN(n23) );
  OAI221_X2 U452 ( .B1(n16400), .B2(n13759), .C1(n24), .C2(n13755), .A(n365), 
        .ZN(n364) );
  NAND2_X2 U454 ( .A1(mem_ExecResult[2]), .A2(n13127), .ZN(n24) );
  OAI221_X2 U457 ( .B1(n16387), .B2(n13759), .C1(n25), .C2(n13755), .A(n367), 
        .ZN(n366) );
  NAND2_X2 U459 ( .A1(mem_ExecResult[3]), .A2(n13127), .ZN(n25) );
  NOR4_X2 U461 ( .A1(n368), .A2(n369), .A3(n120), .A4(n119), .ZN(n324) );
  OAI221_X2 U462 ( .B1(n16196), .B2(n13759), .C1(n13756), .C2(n45), .A(n370), 
        .ZN(n119) );
  NAND2_X2 U464 ( .A1(mem_ExecResult[23]), .A2(n13127), .ZN(n45) );
  OAI221_X2 U466 ( .B1(n16195), .B2(n13759), .C1(n13756), .C2(n44), .A(n371), 
        .ZN(n120) );
  NAND2_X2 U468 ( .A1(mem_ExecResult[22]), .A2(n13127), .ZN(n44) );
  NAND2_X2 U470 ( .A1(n16156), .A2(n16157), .ZN(n369) );
  OAI221_X2 U472 ( .B1(n16193), .B2(n13759), .C1(n13756), .C2(n42), .A(n373), 
        .ZN(n372) );
  NAND2_X2 U474 ( .A1(mem_ExecResult[20]), .A2(n13127), .ZN(n42) );
  OAI221_X2 U477 ( .B1(n16194), .B2(n13759), .C1(n13756), .C2(n43), .A(n375), 
        .ZN(n374) );
  NAND2_X2 U479 ( .A1(mem_ExecResult[21]), .A2(n13127), .ZN(n43) );
  NAND4_X2 U481 ( .A1(n16152), .A2(n16153), .A3(n16154), .A4(n16155), .ZN(n368) );
  OAI221_X2 U483 ( .B1(n16296), .B2(n13759), .C1(n38), .C2(n13755), .A(n377), 
        .ZN(n376) );
  NAND2_X2 U485 ( .A1(mem_ExecResult[16]), .A2(n13127), .ZN(n38) );
  OAI221_X2 U488 ( .B1(n16211), .B2(n13759), .C1(n13756), .C2(n39), .A(n379), 
        .ZN(n378) );
  NAND2_X2 U490 ( .A1(mem_ExecResult[17]), .A2(n13126), .ZN(n39) );
  OAI221_X2 U493 ( .B1(n16210), .B2(n13760), .C1(n13756), .C2(n40), .A(n381), 
        .ZN(n380) );
  NAND2_X2 U495 ( .A1(mem_ExecResult[18]), .A2(n13126), .ZN(n40) );
  OAI221_X2 U498 ( .B1(n16209), .B2(n13760), .C1(n13757), .C2(n41), .A(n383), 
        .ZN(n382) );
  NAND2_X2 U500 ( .A1(mem_ExecResult[19]), .A2(n13126), .ZN(n41) );
  NOR4_X2 U502 ( .A1(n118), .A2(n117), .A3(n116), .A4(n115), .ZN(n323) );
  OAI221_X2 U503 ( .B1(n16178), .B2(n13760), .C1(n13757), .C2(n49), .A(n384), 
        .ZN(n115) );
  NAND2_X2 U505 ( .A1(mem_ExecResult[27]), .A2(n13126), .ZN(n49) );
  OAI221_X2 U507 ( .B1(n16190), .B2(n13760), .C1(n13757), .C2(n48), .A(n385), 
        .ZN(n116) );
  NAND2_X2 U509 ( .A1(mem_ExecResult[26]), .A2(n13126), .ZN(n48) );
  OAI221_X2 U511 ( .B1(n16189), .B2(n13760), .C1(n13757), .C2(n47), .A(n386), 
        .ZN(n117) );
  NAND2_X2 U513 ( .A1(mem_ExecResult[25]), .A2(n13126), .ZN(n47) );
  OAI221_X2 U515 ( .B1(n16197), .B2(n13760), .C1(n13757), .C2(n46), .A(n387), 
        .ZN(n118) );
  NAND2_X2 U517 ( .A1(mem_ExecResult[24]), .A2(n13126), .ZN(n46) );
  NOR4_X2 U519 ( .A1(n114), .A2(n113), .A3(n112), .A4(n111), .ZN(n322) );
  OAI221_X2 U520 ( .B1(n16176), .B2(n13760), .C1(n13757), .C2(n53), .A(n388), 
        .ZN(n111) );
  NAND2_X2 U522 ( .A1(mem_ExecResult[31]), .A2(n13126), .ZN(n53) );
  OAI221_X2 U524 ( .B1(n16177), .B2(n13760), .C1(n13757), .C2(n52), .A(n389), 
        .ZN(n112) );
  NAND2_X2 U526 ( .A1(mem_ExecResult[30]), .A2(n13126), .ZN(n52) );
  OAI221_X2 U528 ( .B1(n16180), .B2(n13760), .C1(n13757), .C2(n51), .A(n390), 
        .ZN(n113) );
  NAND2_X2 U530 ( .A1(mem_ExecResult[29]), .A2(n13126), .ZN(n51) );
  OAI221_X2 U532 ( .B1(n16179), .B2(n13760), .C1(n13757), .C2(n50), .A(n391), 
        .ZN(n114) );
  NAND2_X2 U539 ( .A1(mem_ExecResult[28]), .A2(n13126), .ZN(n50) );
  NAND2_X2 U546 ( .A1(decode_regfile_intregs_9__9_), .A2(n13740), .ZN(n397) );
  NAND2_X2 U548 ( .A1(decode_regfile_intregs_9__8_), .A2(n13742), .ZN(n399) );
  NAND2_X2 U550 ( .A1(decode_regfile_intregs_9__7_), .A2(n13742), .ZN(n401) );
  NAND2_X2 U552 ( .A1(decode_regfile_intregs_9__6_), .A2(n13742), .ZN(n403) );
  NAND2_X2 U554 ( .A1(decode_regfile_intregs_9__5_), .A2(n13742), .ZN(n405) );
  NAND2_X2 U556 ( .A1(decode_regfile_intregs_9__4_), .A2(n13742), .ZN(n407) );
  NAND2_X2 U558 ( .A1(decode_regfile_intregs_9__3_), .A2(n13742), .ZN(n409) );
  NAND2_X2 U560 ( .A1(decode_regfile_intregs_9__31_), .A2(n13742), .ZN(n411)
         );
  NAND2_X2 U562 ( .A1(decode_regfile_intregs_9__30_), .A2(n13741), .ZN(n413)
         );
  NAND2_X2 U564 ( .A1(decode_regfile_intregs_9__2_), .A2(n13741), .ZN(n415) );
  NAND2_X2 U566 ( .A1(decode_regfile_intregs_9__29_), .A2(n13741), .ZN(n417)
         );
  NAND2_X2 U568 ( .A1(decode_regfile_intregs_9__28_), .A2(n13741), .ZN(n419)
         );
  NAND2_X2 U570 ( .A1(decode_regfile_intregs_9__27_), .A2(n13741), .ZN(n421)
         );
  NAND2_X2 U572 ( .A1(decode_regfile_intregs_9__26_), .A2(n13741), .ZN(n423)
         );
  NAND2_X2 U574 ( .A1(decode_regfile_intregs_9__25_), .A2(n13741), .ZN(n425)
         );
  NAND2_X2 U576 ( .A1(decode_regfile_intregs_9__24_), .A2(n13741), .ZN(n427)
         );
  NAND2_X2 U578 ( .A1(decode_regfile_intregs_9__23_), .A2(n13741), .ZN(n429)
         );
  NAND2_X2 U580 ( .A1(decode_regfile_intregs_9__22_), .A2(n13741), .ZN(n431)
         );
  NAND2_X2 U582 ( .A1(decode_regfile_intregs_9__21_), .A2(n13741), .ZN(n433)
         );
  NAND2_X2 U584 ( .A1(decode_regfile_intregs_9__20_), .A2(n13741), .ZN(n435)
         );
  NAND2_X2 U586 ( .A1(decode_regfile_intregs_9__1_), .A2(n13741), .ZN(n437) );
  NAND2_X2 U588 ( .A1(decode_regfile_intregs_9__19_), .A2(n13741), .ZN(n439)
         );
  NAND2_X2 U590 ( .A1(decode_regfile_intregs_9__18_), .A2(n13741), .ZN(n441)
         );
  NAND2_X2 U592 ( .A1(decode_regfile_intregs_9__17_), .A2(n13741), .ZN(n443)
         );
  NAND2_X2 U594 ( .A1(decode_regfile_intregs_9__16_), .A2(n13740), .ZN(n445)
         );
  NAND2_X2 U596 ( .A1(decode_regfile_intregs_9__15_), .A2(n13740), .ZN(n447)
         );
  NAND2_X2 U598 ( .A1(decode_regfile_intregs_9__14_), .A2(n13741), .ZN(n449)
         );
  NAND2_X2 U600 ( .A1(decode_regfile_intregs_9__13_), .A2(n13740), .ZN(n451)
         );
  NAND2_X2 U602 ( .A1(decode_regfile_intregs_9__12_), .A2(n13740), .ZN(n453)
         );
  NAND2_X2 U604 ( .A1(decode_regfile_intregs_9__11_), .A2(n13741), .ZN(n455)
         );
  NAND2_X2 U606 ( .A1(decode_regfile_intregs_9__10_), .A2(n13740), .ZN(n457)
         );
  NAND2_X2 U608 ( .A1(decode_regfile_intregs_9__0_), .A2(n13741), .ZN(n459) );
  NAND2_X2 U611 ( .A1(decode_regfile_intregs_8__9_), .A2(n13642), .ZN(n463) );
  NAND2_X2 U613 ( .A1(decode_regfile_intregs_8__8_), .A2(n13644), .ZN(n464) );
  NAND2_X2 U615 ( .A1(decode_regfile_intregs_8__7_), .A2(n13644), .ZN(n465) );
  NAND2_X2 U617 ( .A1(decode_regfile_intregs_8__6_), .A2(n13644), .ZN(n466) );
  NAND2_X2 U619 ( .A1(decode_regfile_intregs_8__5_), .A2(n13644), .ZN(n467) );
  NAND2_X2 U621 ( .A1(decode_regfile_intregs_8__4_), .A2(n13644), .ZN(n468) );
  NAND2_X2 U623 ( .A1(decode_regfile_intregs_8__3_), .A2(n13644), .ZN(n469) );
  NAND2_X2 U625 ( .A1(decode_regfile_intregs_8__31_), .A2(n13644), .ZN(n470)
         );
  NAND2_X2 U627 ( .A1(decode_regfile_intregs_8__30_), .A2(n13643), .ZN(n471)
         );
  NAND2_X2 U629 ( .A1(decode_regfile_intregs_8__2_), .A2(n13643), .ZN(n472) );
  NAND2_X2 U631 ( .A1(decode_regfile_intregs_8__29_), .A2(n13643), .ZN(n473)
         );
  NAND2_X2 U633 ( .A1(decode_regfile_intregs_8__28_), .A2(n13643), .ZN(n474)
         );
  NAND2_X2 U635 ( .A1(decode_regfile_intregs_8__27_), .A2(n13643), .ZN(n475)
         );
  NAND2_X2 U637 ( .A1(decode_regfile_intregs_8__26_), .A2(n13643), .ZN(n476)
         );
  NAND2_X2 U639 ( .A1(decode_regfile_intregs_8__25_), .A2(n13643), .ZN(n477)
         );
  NAND2_X2 U641 ( .A1(decode_regfile_intregs_8__24_), .A2(n13643), .ZN(n478)
         );
  NAND2_X2 U643 ( .A1(decode_regfile_intregs_8__23_), .A2(n13643), .ZN(n479)
         );
  NAND2_X2 U645 ( .A1(decode_regfile_intregs_8__22_), .A2(n13643), .ZN(n480)
         );
  NAND2_X2 U647 ( .A1(decode_regfile_intregs_8__21_), .A2(n13643), .ZN(n481)
         );
  NAND2_X2 U649 ( .A1(decode_regfile_intregs_8__20_), .A2(n13643), .ZN(n482)
         );
  NAND2_X2 U651 ( .A1(decode_regfile_intregs_8__1_), .A2(n13643), .ZN(n483) );
  NAND2_X2 U653 ( .A1(decode_regfile_intregs_8__19_), .A2(n13643), .ZN(n484)
         );
  NAND2_X2 U655 ( .A1(decode_regfile_intregs_8__18_), .A2(n13643), .ZN(n485)
         );
  NAND2_X2 U657 ( .A1(decode_regfile_intregs_8__17_), .A2(n13643), .ZN(n486)
         );
  NAND2_X2 U659 ( .A1(decode_regfile_intregs_8__16_), .A2(n13642), .ZN(n487)
         );
  NAND2_X2 U661 ( .A1(decode_regfile_intregs_8__15_), .A2(n13642), .ZN(n488)
         );
  NAND2_X2 U663 ( .A1(decode_regfile_intregs_8__14_), .A2(n13643), .ZN(n489)
         );
  NAND2_X2 U665 ( .A1(decode_regfile_intregs_8__13_), .A2(n13642), .ZN(n490)
         );
  NAND2_X2 U667 ( .A1(decode_regfile_intregs_8__12_), .A2(n13642), .ZN(n491)
         );
  NAND2_X2 U669 ( .A1(decode_regfile_intregs_8__11_), .A2(n13643), .ZN(n492)
         );
  NAND2_X2 U671 ( .A1(decode_regfile_intregs_8__10_), .A2(n13642), .ZN(n493)
         );
  NAND2_X2 U673 ( .A1(decode_regfile_intregs_8__0_), .A2(n13643), .ZN(n494) );
  NAND2_X2 U676 ( .A1(decode_regfile_intregs_7__9_), .A2(n13637), .ZN(n497) );
  NAND2_X2 U678 ( .A1(decode_regfile_intregs_7__8_), .A2(n13639), .ZN(n498) );
  NAND2_X2 U680 ( .A1(decode_regfile_intregs_7__7_), .A2(n13639), .ZN(n499) );
  NAND2_X2 U682 ( .A1(decode_regfile_intregs_7__6_), .A2(n13639), .ZN(n500) );
  NAND2_X2 U684 ( .A1(decode_regfile_intregs_7__5_), .A2(n13639), .ZN(n501) );
  NAND2_X2 U686 ( .A1(decode_regfile_intregs_7__4_), .A2(n13639), .ZN(n502) );
  NAND2_X2 U688 ( .A1(decode_regfile_intregs_7__3_), .A2(n13639), .ZN(n503) );
  NAND2_X2 U690 ( .A1(decode_regfile_intregs_7__31_), .A2(n13639), .ZN(n504)
         );
  NAND2_X2 U692 ( .A1(decode_regfile_intregs_7__30_), .A2(n13638), .ZN(n505)
         );
  NAND2_X2 U694 ( .A1(decode_regfile_intregs_7__2_), .A2(n13638), .ZN(n506) );
  NAND2_X2 U696 ( .A1(decode_regfile_intregs_7__29_), .A2(n13638), .ZN(n507)
         );
  NAND2_X2 U698 ( .A1(decode_regfile_intregs_7__28_), .A2(n13638), .ZN(n508)
         );
  NAND2_X2 U700 ( .A1(decode_regfile_intregs_7__27_), .A2(n13638), .ZN(n509)
         );
  NAND2_X2 U702 ( .A1(decode_regfile_intregs_7__26_), .A2(n13638), .ZN(n510)
         );
  NAND2_X2 U704 ( .A1(decode_regfile_intregs_7__25_), .A2(n13638), .ZN(n511)
         );
  NAND2_X2 U706 ( .A1(decode_regfile_intregs_7__24_), .A2(n13638), .ZN(n512)
         );
  NAND2_X2 U708 ( .A1(decode_regfile_intregs_7__23_), .A2(n13638), .ZN(n513)
         );
  NAND2_X2 U710 ( .A1(decode_regfile_intregs_7__22_), .A2(n13638), .ZN(n514)
         );
  NAND2_X2 U712 ( .A1(decode_regfile_intregs_7__21_), .A2(n13638), .ZN(n515)
         );
  NAND2_X2 U714 ( .A1(decode_regfile_intregs_7__20_), .A2(n13638), .ZN(n516)
         );
  NAND2_X2 U716 ( .A1(decode_regfile_intregs_7__1_), .A2(n13638), .ZN(n517) );
  NAND2_X2 U718 ( .A1(decode_regfile_intregs_7__19_), .A2(n13638), .ZN(n518)
         );
  NAND2_X2 U720 ( .A1(decode_regfile_intregs_7__18_), .A2(n13638), .ZN(n519)
         );
  NAND2_X2 U722 ( .A1(decode_regfile_intregs_7__17_), .A2(n13638), .ZN(n520)
         );
  NAND2_X2 U724 ( .A1(decode_regfile_intregs_7__16_), .A2(n13637), .ZN(n521)
         );
  NAND2_X2 U726 ( .A1(decode_regfile_intregs_7__15_), .A2(n13637), .ZN(n522)
         );
  NAND2_X2 U728 ( .A1(decode_regfile_intregs_7__14_), .A2(n13638), .ZN(n523)
         );
  NAND2_X2 U730 ( .A1(decode_regfile_intregs_7__13_), .A2(n13637), .ZN(n524)
         );
  NAND2_X2 U732 ( .A1(decode_regfile_intregs_7__12_), .A2(n13637), .ZN(n525)
         );
  NAND2_X2 U734 ( .A1(decode_regfile_intregs_7__11_), .A2(n13638), .ZN(n526)
         );
  NAND2_X2 U736 ( .A1(decode_regfile_intregs_7__10_), .A2(n13637), .ZN(n527)
         );
  NAND2_X2 U738 ( .A1(decode_regfile_intregs_7__0_), .A2(n13638), .ZN(n528) );
  NAND2_X2 U741 ( .A1(decode_regfile_intregs_6__9_), .A2(n13632), .ZN(n532) );
  NAND2_X2 U743 ( .A1(decode_regfile_intregs_6__8_), .A2(n13634), .ZN(n533) );
  NAND2_X2 U745 ( .A1(decode_regfile_intregs_6__7_), .A2(n13634), .ZN(n534) );
  NAND2_X2 U747 ( .A1(decode_regfile_intregs_6__6_), .A2(n13634), .ZN(n535) );
  NAND2_X2 U749 ( .A1(decode_regfile_intregs_6__5_), .A2(n13634), .ZN(n536) );
  NAND2_X2 U751 ( .A1(decode_regfile_intregs_6__4_), .A2(n13634), .ZN(n537) );
  NAND2_X2 U753 ( .A1(decode_regfile_intregs_6__3_), .A2(n13634), .ZN(n538) );
  NAND2_X2 U755 ( .A1(decode_regfile_intregs_6__31_), .A2(n13634), .ZN(n539)
         );
  NAND2_X2 U757 ( .A1(decode_regfile_intregs_6__30_), .A2(n13633), .ZN(n540)
         );
  NAND2_X2 U759 ( .A1(decode_regfile_intregs_6__2_), .A2(n13633), .ZN(n541) );
  NAND2_X2 U761 ( .A1(decode_regfile_intregs_6__29_), .A2(n13633), .ZN(n542)
         );
  NAND2_X2 U763 ( .A1(decode_regfile_intregs_6__28_), .A2(n13633), .ZN(n543)
         );
  NAND2_X2 U765 ( .A1(decode_regfile_intregs_6__27_), .A2(n13633), .ZN(n544)
         );
  NAND2_X2 U767 ( .A1(decode_regfile_intregs_6__26_), .A2(n13633), .ZN(n545)
         );
  NAND2_X2 U769 ( .A1(decode_regfile_intregs_6__25_), .A2(n13633), .ZN(n546)
         );
  NAND2_X2 U771 ( .A1(decode_regfile_intregs_6__24_), .A2(n13633), .ZN(n547)
         );
  NAND2_X2 U773 ( .A1(decode_regfile_intregs_6__23_), .A2(n13633), .ZN(n548)
         );
  NAND2_X2 U775 ( .A1(decode_regfile_intregs_6__22_), .A2(n13633), .ZN(n549)
         );
  NAND2_X2 U777 ( .A1(decode_regfile_intregs_6__21_), .A2(n13633), .ZN(n550)
         );
  NAND2_X2 U779 ( .A1(decode_regfile_intregs_6__20_), .A2(n13633), .ZN(n551)
         );
  NAND2_X2 U781 ( .A1(decode_regfile_intregs_6__1_), .A2(n13633), .ZN(n552) );
  NAND2_X2 U783 ( .A1(decode_regfile_intregs_6__19_), .A2(n13633), .ZN(n553)
         );
  NAND2_X2 U785 ( .A1(decode_regfile_intregs_6__18_), .A2(n13633), .ZN(n554)
         );
  NAND2_X2 U787 ( .A1(decode_regfile_intregs_6__17_), .A2(n13633), .ZN(n555)
         );
  NAND2_X2 U789 ( .A1(decode_regfile_intregs_6__16_), .A2(n13632), .ZN(n556)
         );
  NAND2_X2 U791 ( .A1(decode_regfile_intregs_6__15_), .A2(n13632), .ZN(n557)
         );
  NAND2_X2 U793 ( .A1(decode_regfile_intregs_6__14_), .A2(n13633), .ZN(n558)
         );
  NAND2_X2 U795 ( .A1(decode_regfile_intregs_6__13_), .A2(n13632), .ZN(n559)
         );
  NAND2_X2 U797 ( .A1(decode_regfile_intregs_6__12_), .A2(n13632), .ZN(n560)
         );
  NAND2_X2 U799 ( .A1(decode_regfile_intregs_6__11_), .A2(n13633), .ZN(n561)
         );
  NAND2_X2 U801 ( .A1(decode_regfile_intregs_6__10_), .A2(n13632), .ZN(n562)
         );
  NAND2_X2 U803 ( .A1(decode_regfile_intregs_6__0_), .A2(n13633), .ZN(n563) );
  NAND2_X2 U806 ( .A1(decode_regfile_intregs_5__9_), .A2(n13627), .ZN(n566) );
  NAND2_X2 U808 ( .A1(decode_regfile_intregs_5__8_), .A2(n13629), .ZN(n567) );
  NAND2_X2 U810 ( .A1(decode_regfile_intregs_5__7_), .A2(n13629), .ZN(n568) );
  NAND2_X2 U812 ( .A1(decode_regfile_intregs_5__6_), .A2(n13629), .ZN(n569) );
  NAND2_X2 U814 ( .A1(decode_regfile_intregs_5__5_), .A2(n13629), .ZN(n570) );
  NAND2_X2 U816 ( .A1(decode_regfile_intregs_5__4_), .A2(n13629), .ZN(n571) );
  NAND2_X2 U818 ( .A1(decode_regfile_intregs_5__3_), .A2(n13629), .ZN(n572) );
  NAND2_X2 U820 ( .A1(decode_regfile_intregs_5__31_), .A2(n13629), .ZN(n573)
         );
  NAND2_X2 U822 ( .A1(decode_regfile_intregs_5__30_), .A2(n13628), .ZN(n574)
         );
  NAND2_X2 U824 ( .A1(decode_regfile_intregs_5__2_), .A2(n13628), .ZN(n575) );
  NAND2_X2 U826 ( .A1(decode_regfile_intregs_5__29_), .A2(n13628), .ZN(n576)
         );
  NAND2_X2 U828 ( .A1(decode_regfile_intregs_5__28_), .A2(n13628), .ZN(n577)
         );
  NAND2_X2 U830 ( .A1(decode_regfile_intregs_5__27_), .A2(n13628), .ZN(n578)
         );
  NAND2_X2 U832 ( .A1(decode_regfile_intregs_5__26_), .A2(n13628), .ZN(n579)
         );
  NAND2_X2 U834 ( .A1(decode_regfile_intregs_5__25_), .A2(n13628), .ZN(n580)
         );
  NAND2_X2 U836 ( .A1(decode_regfile_intregs_5__24_), .A2(n13628), .ZN(n581)
         );
  NAND2_X2 U838 ( .A1(decode_regfile_intregs_5__23_), .A2(n13628), .ZN(n582)
         );
  NAND2_X2 U840 ( .A1(decode_regfile_intregs_5__22_), .A2(n13628), .ZN(n583)
         );
  NAND2_X2 U842 ( .A1(decode_regfile_intregs_5__21_), .A2(n13628), .ZN(n584)
         );
  NAND2_X2 U844 ( .A1(decode_regfile_intregs_5__20_), .A2(n13628), .ZN(n585)
         );
  NAND2_X2 U846 ( .A1(decode_regfile_intregs_5__1_), .A2(n13628), .ZN(n586) );
  NAND2_X2 U848 ( .A1(decode_regfile_intregs_5__19_), .A2(n13628), .ZN(n587)
         );
  NAND2_X2 U850 ( .A1(decode_regfile_intregs_5__18_), .A2(n13628), .ZN(n588)
         );
  NAND2_X2 U852 ( .A1(decode_regfile_intregs_5__17_), .A2(n13628), .ZN(n589)
         );
  NAND2_X2 U854 ( .A1(decode_regfile_intregs_5__16_), .A2(n13627), .ZN(n590)
         );
  NAND2_X2 U856 ( .A1(decode_regfile_intregs_5__15_), .A2(n13627), .ZN(n591)
         );
  NAND2_X2 U858 ( .A1(decode_regfile_intregs_5__14_), .A2(n13628), .ZN(n592)
         );
  NAND2_X2 U860 ( .A1(decode_regfile_intregs_5__13_), .A2(n13627), .ZN(n593)
         );
  NAND2_X2 U862 ( .A1(decode_regfile_intregs_5__12_), .A2(n13627), .ZN(n594)
         );
  NAND2_X2 U864 ( .A1(decode_regfile_intregs_5__11_), .A2(n13628), .ZN(n595)
         );
  NAND2_X2 U866 ( .A1(decode_regfile_intregs_5__10_), .A2(n13627), .ZN(n596)
         );
  NAND2_X2 U868 ( .A1(decode_regfile_intregs_5__0_), .A2(n13628), .ZN(n597) );
  NAND2_X2 U871 ( .A1(decode_regfile_intregs_4__9_), .A2(n13622), .ZN(n599) );
  NAND2_X2 U873 ( .A1(decode_regfile_intregs_4__8_), .A2(n13624), .ZN(n600) );
  NAND2_X2 U875 ( .A1(decode_regfile_intregs_4__7_), .A2(n13624), .ZN(n601) );
  NAND2_X2 U877 ( .A1(decode_regfile_intregs_4__6_), .A2(n13624), .ZN(n602) );
  NAND2_X2 U879 ( .A1(decode_regfile_intregs_4__5_), .A2(n13624), .ZN(n603) );
  NAND2_X2 U881 ( .A1(decode_regfile_intregs_4__4_), .A2(n13624), .ZN(n604) );
  NAND2_X2 U883 ( .A1(decode_regfile_intregs_4__3_), .A2(n13624), .ZN(n605) );
  NAND2_X2 U885 ( .A1(decode_regfile_intregs_4__31_), .A2(n13624), .ZN(n606)
         );
  NAND2_X2 U887 ( .A1(decode_regfile_intregs_4__30_), .A2(n13623), .ZN(n607)
         );
  NAND2_X2 U889 ( .A1(decode_regfile_intregs_4__2_), .A2(n13623), .ZN(n608) );
  NAND2_X2 U891 ( .A1(decode_regfile_intregs_4__29_), .A2(n13623), .ZN(n609)
         );
  NAND2_X2 U893 ( .A1(decode_regfile_intregs_4__28_), .A2(n13623), .ZN(n610)
         );
  NAND2_X2 U895 ( .A1(decode_regfile_intregs_4__27_), .A2(n13623), .ZN(n611)
         );
  NAND2_X2 U897 ( .A1(decode_regfile_intregs_4__26_), .A2(n13623), .ZN(n612)
         );
  NAND2_X2 U899 ( .A1(decode_regfile_intregs_4__25_), .A2(n13623), .ZN(n613)
         );
  NAND2_X2 U901 ( .A1(decode_regfile_intregs_4__24_), .A2(n13623), .ZN(n614)
         );
  NAND2_X2 U903 ( .A1(decode_regfile_intregs_4__23_), .A2(n13623), .ZN(n615)
         );
  NAND2_X2 U905 ( .A1(decode_regfile_intregs_4__22_), .A2(n13623), .ZN(n616)
         );
  NAND2_X2 U907 ( .A1(decode_regfile_intregs_4__21_), .A2(n13623), .ZN(n617)
         );
  NAND2_X2 U909 ( .A1(decode_regfile_intregs_4__20_), .A2(n13623), .ZN(n618)
         );
  NAND2_X2 U911 ( .A1(decode_regfile_intregs_4__1_), .A2(n13623), .ZN(n619) );
  NAND2_X2 U913 ( .A1(decode_regfile_intregs_4__19_), .A2(n13623), .ZN(n620)
         );
  NAND2_X2 U915 ( .A1(decode_regfile_intregs_4__18_), .A2(n13623), .ZN(n621)
         );
  NAND2_X2 U917 ( .A1(decode_regfile_intregs_4__17_), .A2(n13623), .ZN(n622)
         );
  NAND2_X2 U919 ( .A1(decode_regfile_intregs_4__16_), .A2(n13622), .ZN(n623)
         );
  NAND2_X2 U921 ( .A1(decode_regfile_intregs_4__15_), .A2(n13622), .ZN(n624)
         );
  NAND2_X2 U923 ( .A1(decode_regfile_intregs_4__14_), .A2(n13623), .ZN(n625)
         );
  NAND2_X2 U925 ( .A1(decode_regfile_intregs_4__13_), .A2(n13622), .ZN(n626)
         );
  NAND2_X2 U927 ( .A1(decode_regfile_intregs_4__12_), .A2(n13622), .ZN(n627)
         );
  NAND2_X2 U929 ( .A1(decode_regfile_intregs_4__11_), .A2(n13623), .ZN(n628)
         );
  NAND2_X2 U931 ( .A1(decode_regfile_intregs_4__10_), .A2(n13622), .ZN(n629)
         );
  NAND2_X2 U933 ( .A1(decode_regfile_intregs_4__0_), .A2(n13623), .ZN(n630) );
  NAND2_X2 U936 ( .A1(decode_regfile_intregs_3__9_), .A2(n13617), .ZN(n632) );
  NAND2_X2 U938 ( .A1(decode_regfile_intregs_3__8_), .A2(n13619), .ZN(n633) );
  NAND2_X2 U940 ( .A1(decode_regfile_intregs_3__7_), .A2(n13619), .ZN(n634) );
  NAND2_X2 U942 ( .A1(decode_regfile_intregs_3__6_), .A2(n13619), .ZN(n635) );
  NAND2_X2 U944 ( .A1(decode_regfile_intregs_3__5_), .A2(n13619), .ZN(n636) );
  NAND2_X2 U946 ( .A1(decode_regfile_intregs_3__4_), .A2(n13619), .ZN(n637) );
  NAND2_X2 U948 ( .A1(decode_regfile_intregs_3__3_), .A2(n13619), .ZN(n638) );
  NAND2_X2 U950 ( .A1(decode_regfile_intregs_3__31_), .A2(n13619), .ZN(n639)
         );
  NAND2_X2 U952 ( .A1(decode_regfile_intregs_3__30_), .A2(n13618), .ZN(n640)
         );
  NAND2_X2 U954 ( .A1(decode_regfile_intregs_3__2_), .A2(n13618), .ZN(n641) );
  NAND2_X2 U956 ( .A1(decode_regfile_intregs_3__29_), .A2(n13618), .ZN(n642)
         );
  NAND2_X2 U958 ( .A1(decode_regfile_intregs_3__28_), .A2(n13618), .ZN(n643)
         );
  NAND2_X2 U960 ( .A1(decode_regfile_intregs_3__27_), .A2(n13618), .ZN(n644)
         );
  NAND2_X2 U962 ( .A1(decode_regfile_intregs_3__26_), .A2(n13618), .ZN(n645)
         );
  NAND2_X2 U964 ( .A1(decode_regfile_intregs_3__25_), .A2(n13618), .ZN(n646)
         );
  NAND2_X2 U966 ( .A1(decode_regfile_intregs_3__24_), .A2(n13618), .ZN(n647)
         );
  NAND2_X2 U968 ( .A1(decode_regfile_intregs_3__23_), .A2(n13618), .ZN(n648)
         );
  NAND2_X2 U970 ( .A1(decode_regfile_intregs_3__22_), .A2(n13618), .ZN(n649)
         );
  NAND2_X2 U972 ( .A1(decode_regfile_intregs_3__21_), .A2(n13618), .ZN(n650)
         );
  NAND2_X2 U974 ( .A1(decode_regfile_intregs_3__20_), .A2(n13618), .ZN(n651)
         );
  NAND2_X2 U976 ( .A1(decode_regfile_intregs_3__1_), .A2(n13618), .ZN(n652) );
  NAND2_X2 U978 ( .A1(decode_regfile_intregs_3__19_), .A2(n13618), .ZN(n653)
         );
  NAND2_X2 U980 ( .A1(decode_regfile_intregs_3__18_), .A2(n13618), .ZN(n654)
         );
  NAND2_X2 U982 ( .A1(decode_regfile_intregs_3__17_), .A2(n13618), .ZN(n655)
         );
  NAND2_X2 U984 ( .A1(decode_regfile_intregs_3__16_), .A2(n13617), .ZN(n656)
         );
  NAND2_X2 U986 ( .A1(decode_regfile_intregs_3__15_), .A2(n13617), .ZN(n657)
         );
  NAND2_X2 U988 ( .A1(decode_regfile_intregs_3__14_), .A2(n13618), .ZN(n658)
         );
  NAND2_X2 U990 ( .A1(decode_regfile_intregs_3__13_), .A2(n13617), .ZN(n659)
         );
  NAND2_X2 U992 ( .A1(decode_regfile_intregs_3__12_), .A2(n13617), .ZN(n660)
         );
  NAND2_X2 U994 ( .A1(decode_regfile_intregs_3__11_), .A2(n13618), .ZN(n661)
         );
  NAND2_X2 U996 ( .A1(decode_regfile_intregs_3__10_), .A2(n13617), .ZN(n662)
         );
  NAND2_X2 U998 ( .A1(decode_regfile_intregs_3__0_), .A2(n13618), .ZN(n663) );
  NAND2_X2 U1001 ( .A1(decode_regfile_intregs_31__9_), .A2(n13612), .ZN(n666)
         );
  NAND2_X2 U1003 ( .A1(decode_regfile_intregs_31__8_), .A2(n13614), .ZN(n667)
         );
  NAND2_X2 U1005 ( .A1(decode_regfile_intregs_31__7_), .A2(n13614), .ZN(n668)
         );
  NAND2_X2 U1007 ( .A1(decode_regfile_intregs_31__6_), .A2(n13614), .ZN(n669)
         );
  NAND2_X2 U1009 ( .A1(decode_regfile_intregs_31__5_), .A2(n13614), .ZN(n670)
         );
  NAND2_X2 U1011 ( .A1(decode_regfile_intregs_31__4_), .A2(n13614), .ZN(n671)
         );
  NAND2_X2 U1013 ( .A1(decode_regfile_intregs_31__3_), .A2(n13614), .ZN(n672)
         );
  NAND2_X2 U1015 ( .A1(decode_regfile_intregs_31__31_), .A2(n13614), .ZN(n673)
         );
  NAND2_X2 U1017 ( .A1(decode_regfile_intregs_31__30_), .A2(n13613), .ZN(n674)
         );
  NAND2_X2 U1019 ( .A1(decode_regfile_intregs_31__2_), .A2(n13613), .ZN(n675)
         );
  NAND2_X2 U1021 ( .A1(decode_regfile_intregs_31__29_), .A2(n13613), .ZN(n676)
         );
  NAND2_X2 U1023 ( .A1(decode_regfile_intregs_31__28_), .A2(n13613), .ZN(n677)
         );
  NAND2_X2 U1025 ( .A1(decode_regfile_intregs_31__27_), .A2(n13613), .ZN(n678)
         );
  NAND2_X2 U1027 ( .A1(decode_regfile_intregs_31__26_), .A2(n13613), .ZN(n679)
         );
  NAND2_X2 U1029 ( .A1(decode_regfile_intregs_31__25_), .A2(n13613), .ZN(n680)
         );
  NAND2_X2 U1031 ( .A1(decode_regfile_intregs_31__24_), .A2(n13613), .ZN(n681)
         );
  NAND2_X2 U1033 ( .A1(decode_regfile_intregs_31__23_), .A2(n13613), .ZN(n682)
         );
  NAND2_X2 U1035 ( .A1(decode_regfile_intregs_31__22_), .A2(n13613), .ZN(n683)
         );
  NAND2_X2 U1037 ( .A1(decode_regfile_intregs_31__21_), .A2(n13613), .ZN(n684)
         );
  NAND2_X2 U1039 ( .A1(decode_regfile_intregs_31__20_), .A2(n13613), .ZN(n685)
         );
  NAND2_X2 U1041 ( .A1(decode_regfile_intregs_31__1_), .A2(n13613), .ZN(n686)
         );
  NAND2_X2 U1043 ( .A1(decode_regfile_intregs_31__19_), .A2(n13613), .ZN(n687)
         );
  NAND2_X2 U1045 ( .A1(decode_regfile_intregs_31__18_), .A2(n13613), .ZN(n688)
         );
  NAND2_X2 U1047 ( .A1(decode_regfile_intregs_31__17_), .A2(n13613), .ZN(n689)
         );
  NAND2_X2 U1049 ( .A1(decode_regfile_intregs_31__16_), .A2(n13612), .ZN(n690)
         );
  NAND2_X2 U1051 ( .A1(decode_regfile_intregs_31__15_), .A2(n13612), .ZN(n691)
         );
  NAND2_X2 U1053 ( .A1(decode_regfile_intregs_31__14_), .A2(n13613), .ZN(n692)
         );
  NAND2_X2 U1055 ( .A1(decode_regfile_intregs_31__13_), .A2(n13612), .ZN(n693)
         );
  NAND2_X2 U1057 ( .A1(decode_regfile_intregs_31__12_), .A2(n13612), .ZN(n694)
         );
  NAND2_X2 U1059 ( .A1(decode_regfile_intregs_31__11_), .A2(n13613), .ZN(n695)
         );
  NAND2_X2 U1061 ( .A1(decode_regfile_intregs_31__10_), .A2(n13612), .ZN(n696)
         );
  NAND2_X2 U1063 ( .A1(decode_regfile_intregs_31__0_), .A2(n13613), .ZN(n697)
         );
  NAND2_X2 U1066 ( .A1(decode_regfile_intregs_30__9_), .A2(n13607), .ZN(n701)
         );
  NAND2_X2 U1068 ( .A1(decode_regfile_intregs_30__8_), .A2(n13609), .ZN(n702)
         );
  NAND2_X2 U1070 ( .A1(decode_regfile_intregs_30__7_), .A2(n13609), .ZN(n703)
         );
  NAND2_X2 U1072 ( .A1(decode_regfile_intregs_30__6_), .A2(n13609), .ZN(n704)
         );
  NAND2_X2 U1074 ( .A1(decode_regfile_intregs_30__5_), .A2(n13609), .ZN(n705)
         );
  NAND2_X2 U1076 ( .A1(decode_regfile_intregs_30__4_), .A2(n13609), .ZN(n706)
         );
  NAND2_X2 U1078 ( .A1(decode_regfile_intregs_30__3_), .A2(n13609), .ZN(n707)
         );
  NAND2_X2 U1080 ( .A1(decode_regfile_intregs_30__31_), .A2(n13609), .ZN(n708)
         );
  NAND2_X2 U1082 ( .A1(decode_regfile_intregs_30__30_), .A2(n13608), .ZN(n709)
         );
  NAND2_X2 U1084 ( .A1(decode_regfile_intregs_30__2_), .A2(n13608), .ZN(n710)
         );
  NAND2_X2 U1086 ( .A1(decode_regfile_intregs_30__29_), .A2(n13608), .ZN(n711)
         );
  NAND2_X2 U1088 ( .A1(decode_regfile_intregs_30__28_), .A2(n13608), .ZN(n712)
         );
  NAND2_X2 U1090 ( .A1(decode_regfile_intregs_30__27_), .A2(n13608), .ZN(n713)
         );
  NAND2_X2 U1092 ( .A1(decode_regfile_intregs_30__26_), .A2(n13608), .ZN(n714)
         );
  NAND2_X2 U1094 ( .A1(decode_regfile_intregs_30__25_), .A2(n13608), .ZN(n715)
         );
  NAND2_X2 U1096 ( .A1(decode_regfile_intregs_30__24_), .A2(n13608), .ZN(n716)
         );
  NAND2_X2 U1098 ( .A1(decode_regfile_intregs_30__23_), .A2(n13608), .ZN(n717)
         );
  NAND2_X2 U1100 ( .A1(decode_regfile_intregs_30__22_), .A2(n13608), .ZN(n718)
         );
  NAND2_X2 U1102 ( .A1(decode_regfile_intregs_30__21_), .A2(n13608), .ZN(n719)
         );
  NAND2_X2 U1104 ( .A1(decode_regfile_intregs_30__20_), .A2(n13608), .ZN(n720)
         );
  NAND2_X2 U1106 ( .A1(decode_regfile_intregs_30__1_), .A2(n13608), .ZN(n721)
         );
  NAND2_X2 U1108 ( .A1(decode_regfile_intregs_30__19_), .A2(n13608), .ZN(n722)
         );
  NAND2_X2 U1110 ( .A1(decode_regfile_intregs_30__18_), .A2(n13608), .ZN(n723)
         );
  NAND2_X2 U1112 ( .A1(decode_regfile_intregs_30__17_), .A2(n13608), .ZN(n724)
         );
  NAND2_X2 U1114 ( .A1(decode_regfile_intregs_30__16_), .A2(n13607), .ZN(n725)
         );
  NAND2_X2 U1116 ( .A1(decode_regfile_intregs_30__15_), .A2(n13607), .ZN(n726)
         );
  NAND2_X2 U1118 ( .A1(decode_regfile_intregs_30__14_), .A2(n13608), .ZN(n727)
         );
  NAND2_X2 U1120 ( .A1(decode_regfile_intregs_30__13_), .A2(n13607), .ZN(n728)
         );
  NAND2_X2 U1122 ( .A1(decode_regfile_intregs_30__12_), .A2(n13607), .ZN(n729)
         );
  NAND2_X2 U1124 ( .A1(decode_regfile_intregs_30__11_), .A2(n13608), .ZN(n730)
         );
  NAND2_X2 U1126 ( .A1(decode_regfile_intregs_30__10_), .A2(n13607), .ZN(n731)
         );
  NAND2_X2 U1128 ( .A1(decode_regfile_intregs_30__0_), .A2(n13608), .ZN(n732)
         );
  NAND2_X2 U1131 ( .A1(decode_regfile_intregs_2__9_), .A2(n13602), .ZN(n735)
         );
  NAND2_X2 U1133 ( .A1(decode_regfile_intregs_2__8_), .A2(n13604), .ZN(n736)
         );
  NAND2_X2 U1135 ( .A1(decode_regfile_intregs_2__7_), .A2(n13604), .ZN(n737)
         );
  NAND2_X2 U1137 ( .A1(decode_regfile_intregs_2__6_), .A2(n13604), .ZN(n738)
         );
  NAND2_X2 U1139 ( .A1(decode_regfile_intregs_2__5_), .A2(n13604), .ZN(n739)
         );
  NAND2_X2 U1141 ( .A1(decode_regfile_intregs_2__4_), .A2(n13604), .ZN(n740)
         );
  NAND2_X2 U1143 ( .A1(decode_regfile_intregs_2__3_), .A2(n13604), .ZN(n741)
         );
  NAND2_X2 U1145 ( .A1(decode_regfile_intregs_2__31_), .A2(n13604), .ZN(n742)
         );
  NAND2_X2 U1147 ( .A1(decode_regfile_intregs_2__30_), .A2(n13603), .ZN(n743)
         );
  NAND2_X2 U1149 ( .A1(decode_regfile_intregs_2__2_), .A2(n13603), .ZN(n744)
         );
  NAND2_X2 U1151 ( .A1(decode_regfile_intregs_2__29_), .A2(n13603), .ZN(n745)
         );
  NAND2_X2 U1153 ( .A1(decode_regfile_intregs_2__28_), .A2(n13603), .ZN(n746)
         );
  NAND2_X2 U1155 ( .A1(decode_regfile_intregs_2__27_), .A2(n13603), .ZN(n747)
         );
  NAND2_X2 U1157 ( .A1(decode_regfile_intregs_2__26_), .A2(n13603), .ZN(n748)
         );
  NAND2_X2 U1159 ( .A1(decode_regfile_intregs_2__25_), .A2(n13603), .ZN(n749)
         );
  NAND2_X2 U1161 ( .A1(decode_regfile_intregs_2__24_), .A2(n13603), .ZN(n750)
         );
  NAND2_X2 U1163 ( .A1(decode_regfile_intregs_2__23_), .A2(n13603), .ZN(n751)
         );
  NAND2_X2 U1165 ( .A1(decode_regfile_intregs_2__22_), .A2(n13603), .ZN(n752)
         );
  NAND2_X2 U1167 ( .A1(decode_regfile_intregs_2__21_), .A2(n13603), .ZN(n753)
         );
  NAND2_X2 U1169 ( .A1(decode_regfile_intregs_2__20_), .A2(n13603), .ZN(n754)
         );
  NAND2_X2 U1171 ( .A1(decode_regfile_intregs_2__1_), .A2(n13603), .ZN(n755)
         );
  NAND2_X2 U1173 ( .A1(decode_regfile_intregs_2__19_), .A2(n13603), .ZN(n756)
         );
  NAND2_X2 U1175 ( .A1(decode_regfile_intregs_2__18_), .A2(n13603), .ZN(n757)
         );
  NAND2_X2 U1177 ( .A1(decode_regfile_intregs_2__17_), .A2(n13603), .ZN(n758)
         );
  NAND2_X2 U1179 ( .A1(decode_regfile_intregs_2__16_), .A2(n13602), .ZN(n759)
         );
  NAND2_X2 U1181 ( .A1(decode_regfile_intregs_2__15_), .A2(n13602), .ZN(n760)
         );
  NAND2_X2 U1183 ( .A1(decode_regfile_intregs_2__14_), .A2(n13603), .ZN(n761)
         );
  NAND2_X2 U1185 ( .A1(decode_regfile_intregs_2__13_), .A2(n13602), .ZN(n762)
         );
  NAND2_X2 U1187 ( .A1(decode_regfile_intregs_2__12_), .A2(n13602), .ZN(n763)
         );
  NAND2_X2 U1189 ( .A1(decode_regfile_intregs_2__11_), .A2(n13603), .ZN(n764)
         );
  NAND2_X2 U1191 ( .A1(decode_regfile_intregs_2__10_), .A2(n13602), .ZN(n765)
         );
  NAND2_X2 U1193 ( .A1(decode_regfile_intregs_2__0_), .A2(n13603), .ZN(n766)
         );
  NAND2_X2 U1196 ( .A1(decode_regfile_intregs_29__9_), .A2(n13597), .ZN(n768)
         );
  NAND2_X2 U1198 ( .A1(decode_regfile_intregs_29__8_), .A2(n767), .ZN(n769) );
  NAND2_X2 U1200 ( .A1(decode_regfile_intregs_29__7_), .A2(n767), .ZN(n770) );
  NAND2_X2 U1202 ( .A1(decode_regfile_intregs_29__6_), .A2(n767), .ZN(n771) );
  NAND2_X2 U1204 ( .A1(decode_regfile_intregs_29__5_), .A2(n767), .ZN(n772) );
  NAND2_X2 U1206 ( .A1(decode_regfile_intregs_29__4_), .A2(n767), .ZN(n773) );
  NAND2_X2 U1208 ( .A1(decode_regfile_intregs_29__3_), .A2(n767), .ZN(n774) );
  NAND2_X2 U1210 ( .A1(decode_regfile_intregs_29__31_), .A2(n767), .ZN(n775)
         );
  NAND2_X2 U1212 ( .A1(decode_regfile_intregs_29__30_), .A2(n13598), .ZN(n776)
         );
  NAND2_X2 U1214 ( .A1(decode_regfile_intregs_29__2_), .A2(n13598), .ZN(n777)
         );
  NAND2_X2 U1216 ( .A1(decode_regfile_intregs_29__29_), .A2(n13598), .ZN(n778)
         );
  NAND2_X2 U1218 ( .A1(decode_regfile_intregs_29__28_), .A2(n13598), .ZN(n779)
         );
  NAND2_X2 U1220 ( .A1(decode_regfile_intregs_29__27_), .A2(n13598), .ZN(n780)
         );
  NAND2_X2 U1222 ( .A1(decode_regfile_intregs_29__26_), .A2(n13598), .ZN(n781)
         );
  NAND2_X2 U1224 ( .A1(decode_regfile_intregs_29__25_), .A2(n13598), .ZN(n782)
         );
  NAND2_X2 U1226 ( .A1(decode_regfile_intregs_29__24_), .A2(n13598), .ZN(n783)
         );
  NAND2_X2 U1228 ( .A1(decode_regfile_intregs_29__23_), .A2(n13598), .ZN(n784)
         );
  NAND2_X2 U1230 ( .A1(decode_regfile_intregs_29__22_), .A2(n13598), .ZN(n785)
         );
  NAND2_X2 U1232 ( .A1(decode_regfile_intregs_29__21_), .A2(n13598), .ZN(n786)
         );
  NAND2_X2 U1234 ( .A1(decode_regfile_intregs_29__20_), .A2(n13598), .ZN(n787)
         );
  NAND2_X2 U1236 ( .A1(decode_regfile_intregs_29__1_), .A2(n13598), .ZN(n788)
         );
  NAND2_X2 U1238 ( .A1(decode_regfile_intregs_29__19_), .A2(n13598), .ZN(n789)
         );
  NAND2_X2 U1240 ( .A1(decode_regfile_intregs_29__18_), .A2(n13598), .ZN(n790)
         );
  NAND2_X2 U1242 ( .A1(decode_regfile_intregs_29__17_), .A2(n13598), .ZN(n791)
         );
  NAND2_X2 U1244 ( .A1(decode_regfile_intregs_29__16_), .A2(n13597), .ZN(n792)
         );
  NAND2_X2 U1246 ( .A1(decode_regfile_intregs_29__15_), .A2(n13597), .ZN(n793)
         );
  NAND2_X2 U1248 ( .A1(decode_regfile_intregs_29__14_), .A2(n13598), .ZN(n794)
         );
  NAND2_X2 U1250 ( .A1(decode_regfile_intregs_29__13_), .A2(n13597), .ZN(n795)
         );
  NAND2_X2 U1252 ( .A1(decode_regfile_intregs_29__12_), .A2(n13597), .ZN(n796)
         );
  NAND2_X2 U1254 ( .A1(decode_regfile_intregs_29__11_), .A2(n13598), .ZN(n797)
         );
  NAND2_X2 U1256 ( .A1(decode_regfile_intregs_29__10_), .A2(n13597), .ZN(n798)
         );
  NAND2_X2 U1258 ( .A1(decode_regfile_intregs_29__0_), .A2(n13598), .ZN(n799)
         );
  NAND2_X2 U1259 ( .A1(n698), .A2(n800), .ZN(n767) );
  NAND2_X2 U1261 ( .A1(decode_regfile_intregs_28__9_), .A2(n13592), .ZN(n802)
         );
  NAND2_X2 U1263 ( .A1(decode_regfile_intregs_28__8_), .A2(n801), .ZN(n803) );
  NAND2_X2 U1265 ( .A1(decode_regfile_intregs_28__7_), .A2(n801), .ZN(n804) );
  NAND2_X2 U1267 ( .A1(decode_regfile_intregs_28__6_), .A2(n801), .ZN(n805) );
  NAND2_X2 U1269 ( .A1(decode_regfile_intregs_28__5_), .A2(n801), .ZN(n806) );
  NAND2_X2 U1271 ( .A1(decode_regfile_intregs_28__4_), .A2(n801), .ZN(n807) );
  NAND2_X2 U1273 ( .A1(decode_regfile_intregs_28__3_), .A2(n801), .ZN(n808) );
  NAND2_X2 U1275 ( .A1(decode_regfile_intregs_28__31_), .A2(n801), .ZN(n809)
         );
  NAND2_X2 U1277 ( .A1(decode_regfile_intregs_28__30_), .A2(n13593), .ZN(n810)
         );
  NAND2_X2 U1279 ( .A1(decode_regfile_intregs_28__2_), .A2(n13593), .ZN(n811)
         );
  NAND2_X2 U1281 ( .A1(decode_regfile_intregs_28__29_), .A2(n13593), .ZN(n812)
         );
  NAND2_X2 U1283 ( .A1(decode_regfile_intregs_28__28_), .A2(n13593), .ZN(n813)
         );
  NAND2_X2 U1285 ( .A1(decode_regfile_intregs_28__27_), .A2(n13593), .ZN(n814)
         );
  NAND2_X2 U1287 ( .A1(decode_regfile_intregs_28__26_), .A2(n13593), .ZN(n815)
         );
  NAND2_X2 U1289 ( .A1(decode_regfile_intregs_28__25_), .A2(n13593), .ZN(n816)
         );
  NAND2_X2 U1291 ( .A1(decode_regfile_intregs_28__24_), .A2(n13593), .ZN(n817)
         );
  NAND2_X2 U1293 ( .A1(decode_regfile_intregs_28__23_), .A2(n13593), .ZN(n818)
         );
  NAND2_X2 U1295 ( .A1(decode_regfile_intregs_28__22_), .A2(n13593), .ZN(n819)
         );
  NAND2_X2 U1297 ( .A1(decode_regfile_intregs_28__21_), .A2(n13593), .ZN(n820)
         );
  NAND2_X2 U1299 ( .A1(decode_regfile_intregs_28__20_), .A2(n13593), .ZN(n821)
         );
  NAND2_X2 U1301 ( .A1(decode_regfile_intregs_28__1_), .A2(n13593), .ZN(n822)
         );
  NAND2_X2 U1303 ( .A1(decode_regfile_intregs_28__19_), .A2(n13593), .ZN(n823)
         );
  NAND2_X2 U1305 ( .A1(decode_regfile_intregs_28__18_), .A2(n13593), .ZN(n824)
         );
  NAND2_X2 U1307 ( .A1(decode_regfile_intregs_28__17_), .A2(n13593), .ZN(n825)
         );
  NAND2_X2 U1309 ( .A1(decode_regfile_intregs_28__16_), .A2(n13592), .ZN(n826)
         );
  NAND2_X2 U1311 ( .A1(decode_regfile_intregs_28__15_), .A2(n13592), .ZN(n827)
         );
  NAND2_X2 U1313 ( .A1(decode_regfile_intregs_28__14_), .A2(n13593), .ZN(n828)
         );
  NAND2_X2 U1315 ( .A1(decode_regfile_intregs_28__13_), .A2(n13592), .ZN(n829)
         );
  NAND2_X2 U1317 ( .A1(decode_regfile_intregs_28__12_), .A2(n13592), .ZN(n830)
         );
  NAND2_X2 U1319 ( .A1(decode_regfile_intregs_28__11_), .A2(n13593), .ZN(n831)
         );
  NAND2_X2 U1321 ( .A1(decode_regfile_intregs_28__10_), .A2(n13592), .ZN(n832)
         );
  NAND2_X2 U1323 ( .A1(decode_regfile_intregs_28__0_), .A2(n13593), .ZN(n833)
         );
  NAND2_X2 U1324 ( .A1(n698), .A2(n834), .ZN(n801) );
  AND2_X2 U1325 ( .A1(n835), .A2(n836), .ZN(n698) );
  NAND2_X2 U1327 ( .A1(decode_regfile_intregs_27__9_), .A2(n13587), .ZN(n838)
         );
  NAND2_X2 U1329 ( .A1(decode_regfile_intregs_27__8_), .A2(n13589), .ZN(n839)
         );
  NAND2_X2 U1331 ( .A1(decode_regfile_intregs_27__7_), .A2(n13589), .ZN(n840)
         );
  NAND2_X2 U1333 ( .A1(decode_regfile_intregs_27__6_), .A2(n13589), .ZN(n841)
         );
  NAND2_X2 U1335 ( .A1(decode_regfile_intregs_27__5_), .A2(n13589), .ZN(n842)
         );
  NAND2_X2 U1337 ( .A1(decode_regfile_intregs_27__4_), .A2(n13589), .ZN(n843)
         );
  NAND2_X2 U1339 ( .A1(decode_regfile_intregs_27__3_), .A2(n13589), .ZN(n844)
         );
  NAND2_X2 U1341 ( .A1(decode_regfile_intregs_27__31_), .A2(n13589), .ZN(n845)
         );
  NAND2_X2 U1343 ( .A1(decode_regfile_intregs_27__30_), .A2(n13588), .ZN(n846)
         );
  NAND2_X2 U1345 ( .A1(decode_regfile_intregs_27__2_), .A2(n13588), .ZN(n847)
         );
  NAND2_X2 U1347 ( .A1(decode_regfile_intregs_27__29_), .A2(n13588), .ZN(n848)
         );
  NAND2_X2 U1349 ( .A1(decode_regfile_intregs_27__28_), .A2(n13588), .ZN(n849)
         );
  NAND2_X2 U1351 ( .A1(decode_regfile_intregs_27__27_), .A2(n13588), .ZN(n850)
         );
  NAND2_X2 U1353 ( .A1(decode_regfile_intregs_27__26_), .A2(n13588), .ZN(n851)
         );
  NAND2_X2 U1355 ( .A1(decode_regfile_intregs_27__25_), .A2(n13588), .ZN(n852)
         );
  NAND2_X2 U1357 ( .A1(decode_regfile_intregs_27__24_), .A2(n13588), .ZN(n853)
         );
  NAND2_X2 U1359 ( .A1(decode_regfile_intregs_27__23_), .A2(n13588), .ZN(n854)
         );
  NAND2_X2 U1361 ( .A1(decode_regfile_intregs_27__22_), .A2(n13588), .ZN(n855)
         );
  NAND2_X2 U1363 ( .A1(decode_regfile_intregs_27__21_), .A2(n13588), .ZN(n856)
         );
  NAND2_X2 U1365 ( .A1(decode_regfile_intregs_27__20_), .A2(n13588), .ZN(n857)
         );
  NAND2_X2 U1367 ( .A1(decode_regfile_intregs_27__1_), .A2(n13588), .ZN(n858)
         );
  NAND2_X2 U1369 ( .A1(decode_regfile_intregs_27__19_), .A2(n13588), .ZN(n859)
         );
  NAND2_X2 U1371 ( .A1(decode_regfile_intregs_27__18_), .A2(n13588), .ZN(n860)
         );
  NAND2_X2 U1373 ( .A1(decode_regfile_intregs_27__17_), .A2(n13588), .ZN(n861)
         );
  NAND2_X2 U1375 ( .A1(decode_regfile_intregs_27__16_), .A2(n13587), .ZN(n862)
         );
  NAND2_X2 U1377 ( .A1(decode_regfile_intregs_27__15_), .A2(n13587), .ZN(n863)
         );
  NAND2_X2 U1379 ( .A1(decode_regfile_intregs_27__14_), .A2(n13588), .ZN(n864)
         );
  NAND2_X2 U1381 ( .A1(decode_regfile_intregs_27__13_), .A2(n13587), .ZN(n865)
         );
  NAND2_X2 U1383 ( .A1(decode_regfile_intregs_27__12_), .A2(n13587), .ZN(n866)
         );
  NAND2_X2 U1385 ( .A1(decode_regfile_intregs_27__11_), .A2(n13588), .ZN(n867)
         );
  NAND2_X2 U1387 ( .A1(decode_regfile_intregs_27__10_), .A2(n13587), .ZN(n868)
         );
  NAND2_X2 U1389 ( .A1(decode_regfile_intregs_27__0_), .A2(n13588), .ZN(n869)
         );
  NAND2_X2 U1392 ( .A1(decode_regfile_intregs_26__9_), .A2(n13582), .ZN(n872)
         );
  NAND2_X2 U1394 ( .A1(decode_regfile_intregs_26__8_), .A2(n13584), .ZN(n873)
         );
  NAND2_X2 U1396 ( .A1(decode_regfile_intregs_26__7_), .A2(n13584), .ZN(n874)
         );
  NAND2_X2 U1398 ( .A1(decode_regfile_intregs_26__6_), .A2(n13584), .ZN(n875)
         );
  NAND2_X2 U1400 ( .A1(decode_regfile_intregs_26__5_), .A2(n13584), .ZN(n876)
         );
  NAND2_X2 U1402 ( .A1(decode_regfile_intregs_26__4_), .A2(n13584), .ZN(n877)
         );
  NAND2_X2 U1404 ( .A1(decode_regfile_intregs_26__3_), .A2(n13584), .ZN(n878)
         );
  NAND2_X2 U1406 ( .A1(decode_regfile_intregs_26__31_), .A2(n13584), .ZN(n879)
         );
  NAND2_X2 U1408 ( .A1(decode_regfile_intregs_26__30_), .A2(n13583), .ZN(n880)
         );
  NAND2_X2 U1410 ( .A1(decode_regfile_intregs_26__2_), .A2(n13583), .ZN(n881)
         );
  NAND2_X2 U1412 ( .A1(decode_regfile_intregs_26__29_), .A2(n13583), .ZN(n882)
         );
  NAND2_X2 U1414 ( .A1(decode_regfile_intregs_26__28_), .A2(n13583), .ZN(n883)
         );
  NAND2_X2 U1416 ( .A1(decode_regfile_intregs_26__27_), .A2(n13583), .ZN(n884)
         );
  NAND2_X2 U1418 ( .A1(decode_regfile_intregs_26__26_), .A2(n13583), .ZN(n885)
         );
  NAND2_X2 U1420 ( .A1(decode_regfile_intregs_26__25_), .A2(n13583), .ZN(n886)
         );
  NAND2_X2 U1422 ( .A1(decode_regfile_intregs_26__24_), .A2(n13583), .ZN(n887)
         );
  NAND2_X2 U1424 ( .A1(decode_regfile_intregs_26__23_), .A2(n13583), .ZN(n888)
         );
  NAND2_X2 U1426 ( .A1(decode_regfile_intregs_26__22_), .A2(n13583), .ZN(n889)
         );
  NAND2_X2 U1428 ( .A1(decode_regfile_intregs_26__21_), .A2(n13583), .ZN(n890)
         );
  NAND2_X2 U1430 ( .A1(decode_regfile_intregs_26__20_), .A2(n13583), .ZN(n891)
         );
  NAND2_X2 U1432 ( .A1(decode_regfile_intregs_26__1_), .A2(n13583), .ZN(n892)
         );
  NAND2_X2 U1434 ( .A1(decode_regfile_intregs_26__19_), .A2(n13583), .ZN(n893)
         );
  NAND2_X2 U1436 ( .A1(decode_regfile_intregs_26__18_), .A2(n13583), .ZN(n894)
         );
  NAND2_X2 U1438 ( .A1(decode_regfile_intregs_26__17_), .A2(n13583), .ZN(n895)
         );
  NAND2_X2 U1440 ( .A1(decode_regfile_intregs_26__16_), .A2(n13582), .ZN(n896)
         );
  NAND2_X2 U1442 ( .A1(decode_regfile_intregs_26__15_), .A2(n13582), .ZN(n897)
         );
  NAND2_X2 U1444 ( .A1(decode_regfile_intregs_26__14_), .A2(n13583), .ZN(n898)
         );
  NAND2_X2 U1446 ( .A1(decode_regfile_intregs_26__13_), .A2(n13582), .ZN(n899)
         );
  NAND2_X2 U1448 ( .A1(decode_regfile_intregs_26__12_), .A2(n13582), .ZN(n900)
         );
  NAND2_X2 U1450 ( .A1(decode_regfile_intregs_26__11_), .A2(n13583), .ZN(n901)
         );
  NAND2_X2 U1452 ( .A1(decode_regfile_intregs_26__10_), .A2(n13582), .ZN(n902)
         );
  NAND2_X2 U1454 ( .A1(decode_regfile_intregs_26__0_), .A2(n13583), .ZN(n903)
         );
  NAND2_X2 U1457 ( .A1(decode_regfile_intregs_25__9_), .A2(n13577), .ZN(n905)
         );
  NAND2_X2 U1459 ( .A1(decode_regfile_intregs_25__8_), .A2(n904), .ZN(n906) );
  NAND2_X2 U1461 ( .A1(decode_regfile_intregs_25__7_), .A2(n904), .ZN(n907) );
  NAND2_X2 U1463 ( .A1(decode_regfile_intregs_25__6_), .A2(n904), .ZN(n908) );
  NAND2_X2 U1465 ( .A1(decode_regfile_intregs_25__5_), .A2(n904), .ZN(n909) );
  NAND2_X2 U1467 ( .A1(decode_regfile_intregs_25__4_), .A2(n904), .ZN(n910) );
  NAND2_X2 U1469 ( .A1(decode_regfile_intregs_25__3_), .A2(n904), .ZN(n911) );
  NAND2_X2 U1471 ( .A1(decode_regfile_intregs_25__31_), .A2(n904), .ZN(n912)
         );
  NAND2_X2 U1473 ( .A1(decode_regfile_intregs_25__30_), .A2(n13578), .ZN(n913)
         );
  NAND2_X2 U1475 ( .A1(decode_regfile_intregs_25__2_), .A2(n13578), .ZN(n914)
         );
  NAND2_X2 U1477 ( .A1(decode_regfile_intregs_25__29_), .A2(n13578), .ZN(n915)
         );
  NAND2_X2 U1479 ( .A1(decode_regfile_intregs_25__28_), .A2(n13578), .ZN(n916)
         );
  NAND2_X2 U1481 ( .A1(decode_regfile_intregs_25__27_), .A2(n13578), .ZN(n917)
         );
  NAND2_X2 U1483 ( .A1(decode_regfile_intregs_25__26_), .A2(n13578), .ZN(n918)
         );
  NAND2_X2 U1485 ( .A1(decode_regfile_intregs_25__25_), .A2(n13578), .ZN(n919)
         );
  NAND2_X2 U1487 ( .A1(decode_regfile_intregs_25__24_), .A2(n13578), .ZN(n920)
         );
  NAND2_X2 U1489 ( .A1(decode_regfile_intregs_25__23_), .A2(n13578), .ZN(n921)
         );
  NAND2_X2 U1491 ( .A1(decode_regfile_intregs_25__22_), .A2(n13578), .ZN(n922)
         );
  NAND2_X2 U1493 ( .A1(decode_regfile_intregs_25__21_), .A2(n13578), .ZN(n923)
         );
  NAND2_X2 U1495 ( .A1(decode_regfile_intregs_25__20_), .A2(n13578), .ZN(n924)
         );
  NAND2_X2 U1497 ( .A1(decode_regfile_intregs_25__1_), .A2(n13578), .ZN(n925)
         );
  NAND2_X2 U1499 ( .A1(decode_regfile_intregs_25__19_), .A2(n13578), .ZN(n926)
         );
  NAND2_X2 U1501 ( .A1(decode_regfile_intregs_25__18_), .A2(n13578), .ZN(n927)
         );
  NAND2_X2 U1503 ( .A1(decode_regfile_intregs_25__17_), .A2(n13578), .ZN(n928)
         );
  NAND2_X2 U1505 ( .A1(decode_regfile_intregs_25__16_), .A2(n13577), .ZN(n929)
         );
  NAND2_X2 U1507 ( .A1(decode_regfile_intregs_25__15_), .A2(n13577), .ZN(n930)
         );
  NAND2_X2 U1509 ( .A1(decode_regfile_intregs_25__14_), .A2(n13578), .ZN(n931)
         );
  NAND2_X2 U1511 ( .A1(decode_regfile_intregs_25__13_), .A2(n13577), .ZN(n932)
         );
  NAND2_X2 U1513 ( .A1(decode_regfile_intregs_25__12_), .A2(n13577), .ZN(n933)
         );
  NAND2_X2 U1515 ( .A1(decode_regfile_intregs_25__11_), .A2(n13578), .ZN(n934)
         );
  NAND2_X2 U1517 ( .A1(decode_regfile_intregs_25__10_), .A2(n13577), .ZN(n935)
         );
  NAND2_X2 U1519 ( .A1(decode_regfile_intregs_25__0_), .A2(n13578), .ZN(n936)
         );
  NAND2_X2 U1520 ( .A1(n870), .A2(n800), .ZN(n904) );
  NAND2_X2 U1522 ( .A1(decode_regfile_intregs_24__9_), .A2(n13572), .ZN(n938)
         );
  NAND2_X2 U1524 ( .A1(decode_regfile_intregs_24__8_), .A2(n937), .ZN(n939) );
  NAND2_X2 U1526 ( .A1(decode_regfile_intregs_24__7_), .A2(n937), .ZN(n940) );
  NAND2_X2 U1528 ( .A1(decode_regfile_intregs_24__6_), .A2(n937), .ZN(n941) );
  NAND2_X2 U1530 ( .A1(decode_regfile_intregs_24__5_), .A2(n937), .ZN(n942) );
  NAND2_X2 U1532 ( .A1(decode_regfile_intregs_24__4_), .A2(n937), .ZN(n943) );
  NAND2_X2 U1534 ( .A1(decode_regfile_intregs_24__3_), .A2(n937), .ZN(n944) );
  NAND2_X2 U1536 ( .A1(decode_regfile_intregs_24__31_), .A2(n937), .ZN(n945)
         );
  NAND2_X2 U1538 ( .A1(decode_regfile_intregs_24__30_), .A2(n13573), .ZN(n946)
         );
  NAND2_X2 U1540 ( .A1(decode_regfile_intregs_24__2_), .A2(n13573), .ZN(n947)
         );
  NAND2_X2 U1542 ( .A1(decode_regfile_intregs_24__29_), .A2(n13573), .ZN(n948)
         );
  NAND2_X2 U1544 ( .A1(decode_regfile_intregs_24__28_), .A2(n13573), .ZN(n949)
         );
  NAND2_X2 U1546 ( .A1(decode_regfile_intregs_24__27_), .A2(n13573), .ZN(n950)
         );
  NAND2_X2 U1548 ( .A1(decode_regfile_intregs_24__26_), .A2(n13573), .ZN(n951)
         );
  NAND2_X2 U1550 ( .A1(decode_regfile_intregs_24__25_), .A2(n13573), .ZN(n952)
         );
  NAND2_X2 U1552 ( .A1(decode_regfile_intregs_24__24_), .A2(n13573), .ZN(n953)
         );
  NAND2_X2 U1554 ( .A1(decode_regfile_intregs_24__23_), .A2(n13573), .ZN(n954)
         );
  NAND2_X2 U1556 ( .A1(decode_regfile_intregs_24__22_), .A2(n13573), .ZN(n955)
         );
  NAND2_X2 U1558 ( .A1(decode_regfile_intregs_24__21_), .A2(n13573), .ZN(n956)
         );
  NAND2_X2 U1560 ( .A1(decode_regfile_intregs_24__20_), .A2(n13573), .ZN(n957)
         );
  NAND2_X2 U1562 ( .A1(decode_regfile_intregs_24__1_), .A2(n13573), .ZN(n958)
         );
  NAND2_X2 U1564 ( .A1(decode_regfile_intregs_24__19_), .A2(n13573), .ZN(n959)
         );
  NAND2_X2 U1566 ( .A1(decode_regfile_intregs_24__18_), .A2(n13573), .ZN(n960)
         );
  NAND2_X2 U1568 ( .A1(decode_regfile_intregs_24__17_), .A2(n13573), .ZN(n961)
         );
  NAND2_X2 U1570 ( .A1(decode_regfile_intregs_24__16_), .A2(n13572), .ZN(n962)
         );
  NAND2_X2 U1572 ( .A1(decode_regfile_intregs_24__15_), .A2(n13572), .ZN(n963)
         );
  NAND2_X2 U1574 ( .A1(decode_regfile_intregs_24__14_), .A2(n13573), .ZN(n964)
         );
  NAND2_X2 U1576 ( .A1(decode_regfile_intregs_24__13_), .A2(n13572), .ZN(n965)
         );
  NAND2_X2 U1578 ( .A1(decode_regfile_intregs_24__12_), .A2(n13572), .ZN(n966)
         );
  NAND2_X2 U1580 ( .A1(decode_regfile_intregs_24__11_), .A2(n13573), .ZN(n967)
         );
  NAND2_X2 U1582 ( .A1(decode_regfile_intregs_24__10_), .A2(n13572), .ZN(n968)
         );
  NAND2_X2 U1584 ( .A1(decode_regfile_intregs_24__0_), .A2(n13573), .ZN(n969)
         );
  NAND2_X2 U1585 ( .A1(n870), .A2(n834), .ZN(n937) );
  AND2_X2 U1586 ( .A1(n835), .A2(n461), .ZN(n870) );
  NAND2_X2 U1588 ( .A1(decode_regfile_intregs_23__9_), .A2(n13567), .ZN(n971)
         );
  NAND2_X2 U1590 ( .A1(decode_regfile_intregs_23__8_), .A2(n13569), .ZN(n972)
         );
  NAND2_X2 U1592 ( .A1(decode_regfile_intregs_23__7_), .A2(n13569), .ZN(n973)
         );
  NAND2_X2 U1594 ( .A1(decode_regfile_intregs_23__6_), .A2(n13569), .ZN(n974)
         );
  NAND2_X2 U1596 ( .A1(decode_regfile_intregs_23__5_), .A2(n13569), .ZN(n975)
         );
  NAND2_X2 U1598 ( .A1(decode_regfile_intregs_23__4_), .A2(n13569), .ZN(n976)
         );
  NAND2_X2 U1600 ( .A1(decode_regfile_intregs_23__3_), .A2(n13569), .ZN(n977)
         );
  NAND2_X2 U1602 ( .A1(decode_regfile_intregs_23__31_), .A2(n13569), .ZN(n978)
         );
  NAND2_X2 U1604 ( .A1(decode_regfile_intregs_23__30_), .A2(n13568), .ZN(n979)
         );
  NAND2_X2 U1606 ( .A1(decode_regfile_intregs_23__2_), .A2(n13568), .ZN(n980)
         );
  NAND2_X2 U1608 ( .A1(decode_regfile_intregs_23__29_), .A2(n13568), .ZN(n981)
         );
  NAND2_X2 U1610 ( .A1(decode_regfile_intregs_23__28_), .A2(n13568), .ZN(n982)
         );
  NAND2_X2 U1612 ( .A1(decode_regfile_intregs_23__27_), .A2(n13568), .ZN(n983)
         );
  NAND2_X2 U1614 ( .A1(decode_regfile_intregs_23__26_), .A2(n13568), .ZN(n984)
         );
  NAND2_X2 U1616 ( .A1(decode_regfile_intregs_23__25_), .A2(n13568), .ZN(n985)
         );
  NAND2_X2 U1618 ( .A1(decode_regfile_intregs_23__24_), .A2(n13568), .ZN(n986)
         );
  NAND2_X2 U1620 ( .A1(decode_regfile_intregs_23__23_), .A2(n13568), .ZN(n987)
         );
  NAND2_X2 U1622 ( .A1(decode_regfile_intregs_23__22_), .A2(n13568), .ZN(n988)
         );
  NAND2_X2 U1624 ( .A1(decode_regfile_intregs_23__21_), .A2(n13568), .ZN(n989)
         );
  NAND2_X2 U1626 ( .A1(decode_regfile_intregs_23__20_), .A2(n13568), .ZN(n990)
         );
  NAND2_X2 U1628 ( .A1(decode_regfile_intregs_23__1_), .A2(n13568), .ZN(n991)
         );
  NAND2_X2 U1630 ( .A1(decode_regfile_intregs_23__19_), .A2(n13568), .ZN(n992)
         );
  NAND2_X2 U1632 ( .A1(decode_regfile_intregs_23__18_), .A2(n13568), .ZN(n993)
         );
  NAND2_X2 U1634 ( .A1(decode_regfile_intregs_23__17_), .A2(n13568), .ZN(n994)
         );
  NAND2_X2 U1636 ( .A1(decode_regfile_intregs_23__16_), .A2(n13567), .ZN(n995)
         );
  NAND2_X2 U1638 ( .A1(decode_regfile_intregs_23__15_), .A2(n13567), .ZN(n996)
         );
  NAND2_X2 U1640 ( .A1(decode_regfile_intregs_23__14_), .A2(n13568), .ZN(n997)
         );
  NAND2_X2 U1642 ( .A1(decode_regfile_intregs_23__13_), .A2(n13567), .ZN(n998)
         );
  NAND2_X2 U1644 ( .A1(decode_regfile_intregs_23__12_), .A2(n13567), .ZN(n999)
         );
  NAND2_X2 U1646 ( .A1(decode_regfile_intregs_23__11_), .A2(n13568), .ZN(n1000) );
  NAND2_X2 U1648 ( .A1(decode_regfile_intregs_23__10_), .A2(n13567), .ZN(n1001) );
  NAND2_X2 U1650 ( .A1(decode_regfile_intregs_23__0_), .A2(n13568), .ZN(n1002)
         );
  NAND2_X2 U1653 ( .A1(decode_regfile_intregs_22__9_), .A2(n13562), .ZN(n1005)
         );
  NAND2_X2 U1655 ( .A1(decode_regfile_intregs_22__8_), .A2(n13564), .ZN(n1006)
         );
  NAND2_X2 U1657 ( .A1(decode_regfile_intregs_22__7_), .A2(n13564), .ZN(n1007)
         );
  NAND2_X2 U1659 ( .A1(decode_regfile_intregs_22__6_), .A2(n13564), .ZN(n1008)
         );
  NAND2_X2 U1661 ( .A1(decode_regfile_intregs_22__5_), .A2(n13564), .ZN(n1009)
         );
  NAND2_X2 U1663 ( .A1(decode_regfile_intregs_22__4_), .A2(n13564), .ZN(n1010)
         );
  NAND2_X2 U1665 ( .A1(decode_regfile_intregs_22__3_), .A2(n13564), .ZN(n1011)
         );
  NAND2_X2 U1667 ( .A1(decode_regfile_intregs_22__31_), .A2(n13564), .ZN(n1012) );
  NAND2_X2 U1669 ( .A1(decode_regfile_intregs_22__30_), .A2(n13563), .ZN(n1013) );
  NAND2_X2 U1671 ( .A1(decode_regfile_intregs_22__2_), .A2(n13563), .ZN(n1014)
         );
  NAND2_X2 U1673 ( .A1(decode_regfile_intregs_22__29_), .A2(n13563), .ZN(n1015) );
  NAND2_X2 U1675 ( .A1(decode_regfile_intregs_22__28_), .A2(n13563), .ZN(n1016) );
  NAND2_X2 U1677 ( .A1(decode_regfile_intregs_22__27_), .A2(n13563), .ZN(n1017) );
  NAND2_X2 U1679 ( .A1(decode_regfile_intregs_22__26_), .A2(n13563), .ZN(n1018) );
  NAND2_X2 U1681 ( .A1(decode_regfile_intregs_22__25_), .A2(n13563), .ZN(n1019) );
  NAND2_X2 U1683 ( .A1(decode_regfile_intregs_22__24_), .A2(n13563), .ZN(n1020) );
  NAND2_X2 U1685 ( .A1(decode_regfile_intregs_22__23_), .A2(n13563), .ZN(n1021) );
  NAND2_X2 U1687 ( .A1(decode_regfile_intregs_22__22_), .A2(n13563), .ZN(n1022) );
  NAND2_X2 U1689 ( .A1(decode_regfile_intregs_22__21_), .A2(n13563), .ZN(n1023) );
  NAND2_X2 U1691 ( .A1(decode_regfile_intregs_22__20_), .A2(n13563), .ZN(n1024) );
  NAND2_X2 U1693 ( .A1(decode_regfile_intregs_22__1_), .A2(n13563), .ZN(n1025)
         );
  NAND2_X2 U1695 ( .A1(decode_regfile_intregs_22__19_), .A2(n13563), .ZN(n1026) );
  NAND2_X2 U1697 ( .A1(decode_regfile_intregs_22__18_), .A2(n13563), .ZN(n1027) );
  NAND2_X2 U1699 ( .A1(decode_regfile_intregs_22__17_), .A2(n13563), .ZN(n1028) );
  NAND2_X2 U1701 ( .A1(decode_regfile_intregs_22__16_), .A2(n13562), .ZN(n1029) );
  NAND2_X2 U1703 ( .A1(decode_regfile_intregs_22__15_), .A2(n13562), .ZN(n1030) );
  NAND2_X2 U1705 ( .A1(decode_regfile_intregs_22__14_), .A2(n13563), .ZN(n1031) );
  NAND2_X2 U1707 ( .A1(decode_regfile_intregs_22__13_), .A2(n13562), .ZN(n1032) );
  NAND2_X2 U1709 ( .A1(decode_regfile_intregs_22__12_), .A2(n13562), .ZN(n1033) );
  NAND2_X2 U1711 ( .A1(decode_regfile_intregs_22__11_), .A2(n13563), .ZN(n1034) );
  NAND2_X2 U1713 ( .A1(decode_regfile_intregs_22__10_), .A2(n13562), .ZN(n1035) );
  NAND2_X2 U1715 ( .A1(decode_regfile_intregs_22__0_), .A2(n13563), .ZN(n1036)
         );
  NAND2_X2 U1718 ( .A1(decode_regfile_intregs_21__9_), .A2(n13557), .ZN(n1038)
         );
  NAND2_X2 U1720 ( .A1(decode_regfile_intregs_21__8_), .A2(n1037), .ZN(n1039)
         );
  NAND2_X2 U1722 ( .A1(decode_regfile_intregs_21__7_), .A2(n1037), .ZN(n1040)
         );
  NAND2_X2 U1724 ( .A1(decode_regfile_intregs_21__6_), .A2(n1037), .ZN(n1041)
         );
  NAND2_X2 U1726 ( .A1(decode_regfile_intregs_21__5_), .A2(n1037), .ZN(n1042)
         );
  NAND2_X2 U1728 ( .A1(decode_regfile_intregs_21__4_), .A2(n1037), .ZN(n1043)
         );
  NAND2_X2 U1730 ( .A1(decode_regfile_intregs_21__3_), .A2(n1037), .ZN(n1044)
         );
  NAND2_X2 U1732 ( .A1(decode_regfile_intregs_21__31_), .A2(n1037), .ZN(n1045)
         );
  NAND2_X2 U1734 ( .A1(decode_regfile_intregs_21__30_), .A2(n13558), .ZN(n1046) );
  NAND2_X2 U1736 ( .A1(decode_regfile_intregs_21__2_), .A2(n13558), .ZN(n1047)
         );
  NAND2_X2 U1738 ( .A1(decode_regfile_intregs_21__29_), .A2(n13558), .ZN(n1048) );
  NAND2_X2 U1740 ( .A1(decode_regfile_intregs_21__28_), .A2(n13558), .ZN(n1049) );
  NAND2_X2 U1742 ( .A1(decode_regfile_intregs_21__27_), .A2(n13558), .ZN(n1050) );
  NAND2_X2 U1744 ( .A1(decode_regfile_intregs_21__26_), .A2(n13558), .ZN(n1051) );
  NAND2_X2 U1746 ( .A1(decode_regfile_intregs_21__25_), .A2(n13558), .ZN(n1052) );
  NAND2_X2 U1748 ( .A1(decode_regfile_intregs_21__24_), .A2(n13558), .ZN(n1053) );
  NAND2_X2 U1750 ( .A1(decode_regfile_intregs_21__23_), .A2(n13558), .ZN(n1054) );
  NAND2_X2 U1752 ( .A1(decode_regfile_intregs_21__22_), .A2(n13558), .ZN(n1055) );
  NAND2_X2 U1754 ( .A1(decode_regfile_intregs_21__21_), .A2(n13558), .ZN(n1056) );
  NAND2_X2 U1756 ( .A1(decode_regfile_intregs_21__20_), .A2(n13558), .ZN(n1057) );
  NAND2_X2 U1758 ( .A1(decode_regfile_intregs_21__1_), .A2(n13558), .ZN(n1058)
         );
  NAND2_X2 U1760 ( .A1(decode_regfile_intregs_21__19_), .A2(n13558), .ZN(n1059) );
  NAND2_X2 U1762 ( .A1(decode_regfile_intregs_21__18_), .A2(n13558), .ZN(n1060) );
  NAND2_X2 U1764 ( .A1(decode_regfile_intregs_21__17_), .A2(n13558), .ZN(n1061) );
  NAND2_X2 U1766 ( .A1(decode_regfile_intregs_21__16_), .A2(n13557), .ZN(n1062) );
  NAND2_X2 U1768 ( .A1(decode_regfile_intregs_21__15_), .A2(n13557), .ZN(n1063) );
  NAND2_X2 U1770 ( .A1(decode_regfile_intregs_21__14_), .A2(n13558), .ZN(n1064) );
  NAND2_X2 U1772 ( .A1(decode_regfile_intregs_21__13_), .A2(n13557), .ZN(n1065) );
  NAND2_X2 U1774 ( .A1(decode_regfile_intregs_21__12_), .A2(n13557), .ZN(n1066) );
  NAND2_X2 U1776 ( .A1(decode_regfile_intregs_21__11_), .A2(n13558), .ZN(n1067) );
  NAND2_X2 U1778 ( .A1(decode_regfile_intregs_21__10_), .A2(n13557), .ZN(n1068) );
  NAND2_X2 U1780 ( .A1(decode_regfile_intregs_21__0_), .A2(n13558), .ZN(n1069)
         );
  NAND2_X2 U1781 ( .A1(n1003), .A2(n800), .ZN(n1037) );
  NAND2_X2 U1783 ( .A1(decode_regfile_intregs_20__9_), .A2(n13552), .ZN(n1071)
         );
  NAND2_X2 U1785 ( .A1(decode_regfile_intregs_20__8_), .A2(n1070), .ZN(n1072)
         );
  NAND2_X2 U1787 ( .A1(decode_regfile_intregs_20__7_), .A2(n1070), .ZN(n1073)
         );
  NAND2_X2 U1789 ( .A1(decode_regfile_intregs_20__6_), .A2(n1070), .ZN(n1074)
         );
  NAND2_X2 U1791 ( .A1(decode_regfile_intregs_20__5_), .A2(n1070), .ZN(n1075)
         );
  NAND2_X2 U1793 ( .A1(decode_regfile_intregs_20__4_), .A2(n1070), .ZN(n1076)
         );
  NAND2_X2 U1795 ( .A1(decode_regfile_intregs_20__3_), .A2(n1070), .ZN(n1077)
         );
  NAND2_X2 U1797 ( .A1(decode_regfile_intregs_20__31_), .A2(n1070), .ZN(n1078)
         );
  NAND2_X2 U1799 ( .A1(decode_regfile_intregs_20__30_), .A2(n13553), .ZN(n1079) );
  NAND2_X2 U1801 ( .A1(decode_regfile_intregs_20__2_), .A2(n13553), .ZN(n1080)
         );
  NAND2_X2 U1803 ( .A1(decode_regfile_intregs_20__29_), .A2(n13553), .ZN(n1081) );
  NAND2_X2 U1805 ( .A1(decode_regfile_intregs_20__28_), .A2(n13553), .ZN(n1082) );
  NAND2_X2 U1807 ( .A1(decode_regfile_intregs_20__27_), .A2(n13553), .ZN(n1083) );
  NAND2_X2 U1809 ( .A1(decode_regfile_intregs_20__26_), .A2(n13553), .ZN(n1084) );
  NAND2_X2 U1811 ( .A1(decode_regfile_intregs_20__25_), .A2(n13553), .ZN(n1085) );
  NAND2_X2 U1813 ( .A1(decode_regfile_intregs_20__24_), .A2(n13553), .ZN(n1086) );
  NAND2_X2 U1815 ( .A1(decode_regfile_intregs_20__23_), .A2(n13553), .ZN(n1087) );
  NAND2_X2 U1817 ( .A1(decode_regfile_intregs_20__22_), .A2(n13553), .ZN(n1088) );
  NAND2_X2 U1819 ( .A1(decode_regfile_intregs_20__21_), .A2(n13553), .ZN(n1089) );
  NAND2_X2 U1821 ( .A1(decode_regfile_intregs_20__20_), .A2(n13553), .ZN(n1090) );
  NAND2_X2 U1823 ( .A1(decode_regfile_intregs_20__1_), .A2(n13553), .ZN(n1091)
         );
  NAND2_X2 U1825 ( .A1(decode_regfile_intregs_20__19_), .A2(n13553), .ZN(n1092) );
  NAND2_X2 U1827 ( .A1(decode_regfile_intregs_20__18_), .A2(n13553), .ZN(n1093) );
  NAND2_X2 U1829 ( .A1(decode_regfile_intregs_20__17_), .A2(n13553), .ZN(n1094) );
  NAND2_X2 U1831 ( .A1(decode_regfile_intregs_20__16_), .A2(n13552), .ZN(n1095) );
  NAND2_X2 U1833 ( .A1(decode_regfile_intregs_20__15_), .A2(n13552), .ZN(n1096) );
  NAND2_X2 U1835 ( .A1(decode_regfile_intregs_20__14_), .A2(n13553), .ZN(n1097) );
  NAND2_X2 U1837 ( .A1(decode_regfile_intregs_20__13_), .A2(n13552), .ZN(n1098) );
  NAND2_X2 U1839 ( .A1(decode_regfile_intregs_20__12_), .A2(n13552), .ZN(n1099) );
  NAND2_X2 U1841 ( .A1(decode_regfile_intregs_20__11_), .A2(n13553), .ZN(n1100) );
  NAND2_X2 U1843 ( .A1(decode_regfile_intregs_20__10_), .A2(n13552), .ZN(n1101) );
  NAND2_X2 U1845 ( .A1(decode_regfile_intregs_20__0_), .A2(n13553), .ZN(n1102)
         );
  NAND2_X2 U1846 ( .A1(n1003), .A2(n834), .ZN(n1070) );
  AND2_X2 U1847 ( .A1(n835), .A2(n530), .ZN(n1003) );
  NAND2_X2 U1849 ( .A1(decode_regfile_intregs_1__9_), .A2(n13547), .ZN(n1104)
         );
  NAND2_X2 U1851 ( .A1(decode_regfile_intregs_1__8_), .A2(n13549), .ZN(n1105)
         );
  NAND2_X2 U1853 ( .A1(decode_regfile_intregs_1__7_), .A2(n13549), .ZN(n1106)
         );
  NAND2_X2 U1855 ( .A1(decode_regfile_intregs_1__6_), .A2(n13549), .ZN(n1107)
         );
  NAND2_X2 U1857 ( .A1(decode_regfile_intregs_1__5_), .A2(n13549), .ZN(n1108)
         );
  NAND2_X2 U1859 ( .A1(decode_regfile_intregs_1__4_), .A2(n13549), .ZN(n1109)
         );
  NAND2_X2 U1861 ( .A1(decode_regfile_intregs_1__3_), .A2(n13549), .ZN(n1110)
         );
  NAND2_X2 U1863 ( .A1(decode_regfile_intregs_1__31_), .A2(n13549), .ZN(n1111)
         );
  NAND2_X2 U1865 ( .A1(decode_regfile_intregs_1__30_), .A2(n13548), .ZN(n1112)
         );
  NAND2_X2 U1867 ( .A1(decode_regfile_intregs_1__2_), .A2(n13548), .ZN(n1113)
         );
  NAND2_X2 U1869 ( .A1(decode_regfile_intregs_1__29_), .A2(n13548), .ZN(n1114)
         );
  NAND2_X2 U1871 ( .A1(decode_regfile_intregs_1__28_), .A2(n13548), .ZN(n1115)
         );
  NAND2_X2 U1873 ( .A1(decode_regfile_intregs_1__27_), .A2(n13548), .ZN(n1116)
         );
  NAND2_X2 U1875 ( .A1(decode_regfile_intregs_1__26_), .A2(n13548), .ZN(n1117)
         );
  NAND2_X2 U1877 ( .A1(decode_regfile_intregs_1__25_), .A2(n13548), .ZN(n1118)
         );
  NAND2_X2 U1879 ( .A1(decode_regfile_intregs_1__24_), .A2(n13548), .ZN(n1119)
         );
  NAND2_X2 U1881 ( .A1(decode_regfile_intregs_1__23_), .A2(n13548), .ZN(n1120)
         );
  NAND2_X2 U1883 ( .A1(decode_regfile_intregs_1__22_), .A2(n13548), .ZN(n1121)
         );
  NAND2_X2 U1885 ( .A1(decode_regfile_intregs_1__21_), .A2(n13548), .ZN(n1122)
         );
  NAND2_X2 U1887 ( .A1(decode_regfile_intregs_1__20_), .A2(n13548), .ZN(n1123)
         );
  NAND2_X2 U1889 ( .A1(decode_regfile_intregs_1__1_), .A2(n13548), .ZN(n1124)
         );
  NAND2_X2 U1891 ( .A1(decode_regfile_intregs_1__19_), .A2(n13548), .ZN(n1125)
         );
  NAND2_X2 U1893 ( .A1(decode_regfile_intregs_1__18_), .A2(n13548), .ZN(n1126)
         );
  NAND2_X2 U1895 ( .A1(decode_regfile_intregs_1__17_), .A2(n13548), .ZN(n1127)
         );
  NAND2_X2 U1897 ( .A1(decode_regfile_intregs_1__16_), .A2(n13547), .ZN(n1128)
         );
  NAND2_X2 U1899 ( .A1(decode_regfile_intregs_1__15_), .A2(n13547), .ZN(n1129)
         );
  NAND2_X2 U1901 ( .A1(decode_regfile_intregs_1__14_), .A2(n13548), .ZN(n1130)
         );
  NAND2_X2 U1903 ( .A1(decode_regfile_intregs_1__13_), .A2(n13547), .ZN(n1131)
         );
  NAND2_X2 U1905 ( .A1(decode_regfile_intregs_1__12_), .A2(n13547), .ZN(n1132)
         );
  NAND2_X2 U1907 ( .A1(decode_regfile_intregs_1__11_), .A2(n13548), .ZN(n1133)
         );
  NAND2_X2 U1909 ( .A1(decode_regfile_intregs_1__10_), .A2(n13547), .ZN(n1134)
         );
  NAND2_X2 U1911 ( .A1(decode_regfile_intregs_1__0_), .A2(n13548), .ZN(n1135)
         );
  NAND2_X2 U1914 ( .A1(decode_regfile_intregs_19__9_), .A2(n13542), .ZN(n1137)
         );
  NAND2_X2 U1916 ( .A1(decode_regfile_intregs_19__8_), .A2(n13544), .ZN(n1138)
         );
  NAND2_X2 U1918 ( .A1(decode_regfile_intregs_19__7_), .A2(n13544), .ZN(n1139)
         );
  NAND2_X2 U1920 ( .A1(decode_regfile_intregs_19__6_), .A2(n13544), .ZN(n1140)
         );
  NAND2_X2 U1922 ( .A1(decode_regfile_intregs_19__5_), .A2(n13544), .ZN(n1141)
         );
  NAND2_X2 U1924 ( .A1(decode_regfile_intregs_19__4_), .A2(n13544), .ZN(n1142)
         );
  NAND2_X2 U1926 ( .A1(decode_regfile_intregs_19__3_), .A2(n13544), .ZN(n1143)
         );
  NAND2_X2 U1928 ( .A1(decode_regfile_intregs_19__31_), .A2(n13544), .ZN(n1144) );
  NAND2_X2 U1930 ( .A1(decode_regfile_intregs_19__30_), .A2(n13543), .ZN(n1145) );
  NAND2_X2 U1932 ( .A1(decode_regfile_intregs_19__2_), .A2(n13543), .ZN(n1146)
         );
  NAND2_X2 U1934 ( .A1(decode_regfile_intregs_19__29_), .A2(n13543), .ZN(n1147) );
  NAND2_X2 U1936 ( .A1(decode_regfile_intregs_19__28_), .A2(n13543), .ZN(n1148) );
  NAND2_X2 U1938 ( .A1(decode_regfile_intregs_19__27_), .A2(n13543), .ZN(n1149) );
  NAND2_X2 U1940 ( .A1(decode_regfile_intregs_19__26_), .A2(n13543), .ZN(n1150) );
  NAND2_X2 U1942 ( .A1(decode_regfile_intregs_19__25_), .A2(n13543), .ZN(n1151) );
  NAND2_X2 U1944 ( .A1(decode_regfile_intregs_19__24_), .A2(n13543), .ZN(n1152) );
  NAND2_X2 U1946 ( .A1(decode_regfile_intregs_19__23_), .A2(n13543), .ZN(n1153) );
  NAND2_X2 U1948 ( .A1(decode_regfile_intregs_19__22_), .A2(n13543), .ZN(n1154) );
  NAND2_X2 U1950 ( .A1(decode_regfile_intregs_19__21_), .A2(n13543), .ZN(n1155) );
  NAND2_X2 U1952 ( .A1(decode_regfile_intregs_19__20_), .A2(n13543), .ZN(n1156) );
  NAND2_X2 U1954 ( .A1(decode_regfile_intregs_19__1_), .A2(n13543), .ZN(n1157)
         );
  NAND2_X2 U1956 ( .A1(decode_regfile_intregs_19__19_), .A2(n13543), .ZN(n1158) );
  NAND2_X2 U1958 ( .A1(decode_regfile_intregs_19__18_), .A2(n13543), .ZN(n1159) );
  NAND2_X2 U1960 ( .A1(decode_regfile_intregs_19__17_), .A2(n13543), .ZN(n1160) );
  NAND2_X2 U1962 ( .A1(decode_regfile_intregs_19__16_), .A2(n13542), .ZN(n1161) );
  NAND2_X2 U1964 ( .A1(decode_regfile_intregs_19__15_), .A2(n13542), .ZN(n1162) );
  NAND2_X2 U1966 ( .A1(decode_regfile_intregs_19__14_), .A2(n13543), .ZN(n1163) );
  NAND2_X2 U1968 ( .A1(decode_regfile_intregs_19__13_), .A2(n13542), .ZN(n1164) );
  NAND2_X2 U1970 ( .A1(decode_regfile_intregs_19__12_), .A2(n13542), .ZN(n1165) );
  NAND2_X2 U1972 ( .A1(decode_regfile_intregs_19__11_), .A2(n13543), .ZN(n1166) );
  NAND2_X2 U1974 ( .A1(decode_regfile_intregs_19__10_), .A2(n13542), .ZN(n1167) );
  NAND2_X2 U1976 ( .A1(decode_regfile_intregs_19__0_), .A2(n13543), .ZN(n1168)
         );
  NAND2_X2 U1979 ( .A1(decode_regfile_intregs_18__9_), .A2(n13537), .ZN(n1171)
         );
  NAND2_X2 U1981 ( .A1(decode_regfile_intregs_18__8_), .A2(n13539), .ZN(n1172)
         );
  NAND2_X2 U1983 ( .A1(decode_regfile_intregs_18__7_), .A2(n13539), .ZN(n1173)
         );
  NAND2_X2 U1985 ( .A1(decode_regfile_intregs_18__6_), .A2(n13539), .ZN(n1174)
         );
  NAND2_X2 U1987 ( .A1(decode_regfile_intregs_18__5_), .A2(n13539), .ZN(n1175)
         );
  NAND2_X2 U1989 ( .A1(decode_regfile_intregs_18__4_), .A2(n13539), .ZN(n1176)
         );
  NAND2_X2 U1991 ( .A1(decode_regfile_intregs_18__3_), .A2(n13539), .ZN(n1177)
         );
  NAND2_X2 U1993 ( .A1(decode_regfile_intregs_18__31_), .A2(n13539), .ZN(n1178) );
  NAND2_X2 U1995 ( .A1(decode_regfile_intregs_18__30_), .A2(n13538), .ZN(n1179) );
  NAND2_X2 U1997 ( .A1(decode_regfile_intregs_18__2_), .A2(n13538), .ZN(n1180)
         );
  NAND2_X2 U1999 ( .A1(decode_regfile_intregs_18__29_), .A2(n13538), .ZN(n1181) );
  NAND2_X2 U2001 ( .A1(decode_regfile_intregs_18__28_), .A2(n13538), .ZN(n1182) );
  NAND2_X2 U2003 ( .A1(decode_regfile_intregs_18__27_), .A2(n13538), .ZN(n1183) );
  NAND2_X2 U2005 ( .A1(decode_regfile_intregs_18__26_), .A2(n13538), .ZN(n1184) );
  NAND2_X2 U2007 ( .A1(decode_regfile_intregs_18__25_), .A2(n13538), .ZN(n1185) );
  NAND2_X2 U2009 ( .A1(decode_regfile_intregs_18__24_), .A2(n13538), .ZN(n1186) );
  NAND2_X2 U2011 ( .A1(decode_regfile_intregs_18__23_), .A2(n13538), .ZN(n1187) );
  NAND2_X2 U2013 ( .A1(decode_regfile_intregs_18__22_), .A2(n13538), .ZN(n1188) );
  NAND2_X2 U2015 ( .A1(decode_regfile_intregs_18__21_), .A2(n13538), .ZN(n1189) );
  NAND2_X2 U2017 ( .A1(decode_regfile_intregs_18__20_), .A2(n13538), .ZN(n1190) );
  NAND2_X2 U2019 ( .A1(decode_regfile_intregs_18__1_), .A2(n13538), .ZN(n1191)
         );
  NAND2_X2 U2021 ( .A1(decode_regfile_intregs_18__19_), .A2(n13538), .ZN(n1192) );
  NAND2_X2 U2023 ( .A1(decode_regfile_intregs_18__18_), .A2(n13538), .ZN(n1193) );
  NAND2_X2 U2025 ( .A1(decode_regfile_intregs_18__17_), .A2(n13538), .ZN(n1194) );
  NAND2_X2 U2027 ( .A1(decode_regfile_intregs_18__16_), .A2(n13537), .ZN(n1195) );
  NAND2_X2 U2029 ( .A1(decode_regfile_intregs_18__15_), .A2(n13537), .ZN(n1196) );
  NAND2_X2 U2031 ( .A1(decode_regfile_intregs_18__14_), .A2(n13538), .ZN(n1197) );
  NAND2_X2 U2033 ( .A1(decode_regfile_intregs_18__13_), .A2(n13537), .ZN(n1198) );
  NAND2_X2 U2035 ( .A1(decode_regfile_intregs_18__12_), .A2(n13537), .ZN(n1199) );
  NAND2_X2 U2037 ( .A1(decode_regfile_intregs_18__11_), .A2(n13538), .ZN(n1200) );
  NAND2_X2 U2039 ( .A1(decode_regfile_intregs_18__10_), .A2(n13537), .ZN(n1201) );
  NAND2_X2 U2041 ( .A1(decode_regfile_intregs_18__0_), .A2(n13538), .ZN(n1202)
         );
  NAND2_X2 U2044 ( .A1(decode_regfile_intregs_17__9_), .A2(n13532), .ZN(n1204)
         );
  NAND2_X2 U2046 ( .A1(decode_regfile_intregs_17__8_), .A2(n1203), .ZN(n1205)
         );
  NAND2_X2 U2048 ( .A1(decode_regfile_intregs_17__7_), .A2(n1203), .ZN(n1206)
         );
  NAND2_X2 U2050 ( .A1(decode_regfile_intregs_17__6_), .A2(n1203), .ZN(n1207)
         );
  NAND2_X2 U2052 ( .A1(decode_regfile_intregs_17__5_), .A2(n1203), .ZN(n1208)
         );
  NAND2_X2 U2054 ( .A1(decode_regfile_intregs_17__4_), .A2(n1203), .ZN(n1209)
         );
  NAND2_X2 U2056 ( .A1(decode_regfile_intregs_17__3_), .A2(n1203), .ZN(n1210)
         );
  NAND2_X2 U2058 ( .A1(decode_regfile_intregs_17__31_), .A2(n1203), .ZN(n1211)
         );
  NAND2_X2 U2060 ( .A1(decode_regfile_intregs_17__30_), .A2(n13533), .ZN(n1212) );
  NAND2_X2 U2062 ( .A1(decode_regfile_intregs_17__2_), .A2(n13533), .ZN(n1213)
         );
  NAND2_X2 U2064 ( .A1(decode_regfile_intregs_17__29_), .A2(n13533), .ZN(n1214) );
  NAND2_X2 U2066 ( .A1(decode_regfile_intregs_17__28_), .A2(n13533), .ZN(n1215) );
  NAND2_X2 U2068 ( .A1(decode_regfile_intregs_17__27_), .A2(n13533), .ZN(n1216) );
  NAND2_X2 U2070 ( .A1(decode_regfile_intregs_17__26_), .A2(n13533), .ZN(n1217) );
  NAND2_X2 U2072 ( .A1(decode_regfile_intregs_17__25_), .A2(n13533), .ZN(n1218) );
  NAND2_X2 U2074 ( .A1(decode_regfile_intregs_17__24_), .A2(n13533), .ZN(n1219) );
  NAND2_X2 U2076 ( .A1(decode_regfile_intregs_17__23_), .A2(n13533), .ZN(n1220) );
  NAND2_X2 U2078 ( .A1(decode_regfile_intregs_17__22_), .A2(n13533), .ZN(n1221) );
  NAND2_X2 U2080 ( .A1(decode_regfile_intregs_17__21_), .A2(n13533), .ZN(n1222) );
  NAND2_X2 U2082 ( .A1(decode_regfile_intregs_17__20_), .A2(n13533), .ZN(n1223) );
  NAND2_X2 U2084 ( .A1(decode_regfile_intregs_17__1_), .A2(n13533), .ZN(n1224)
         );
  NAND2_X2 U2086 ( .A1(decode_regfile_intregs_17__19_), .A2(n13533), .ZN(n1225) );
  NAND2_X2 U2088 ( .A1(decode_regfile_intregs_17__18_), .A2(n13533), .ZN(n1226) );
  NAND2_X2 U2090 ( .A1(decode_regfile_intregs_17__17_), .A2(n13533), .ZN(n1227) );
  NAND2_X2 U2092 ( .A1(decode_regfile_intregs_17__16_), .A2(n13532), .ZN(n1228) );
  NAND2_X2 U2094 ( .A1(decode_regfile_intregs_17__15_), .A2(n13532), .ZN(n1229) );
  NAND2_X2 U2096 ( .A1(decode_regfile_intregs_17__14_), .A2(n13533), .ZN(n1230) );
  NAND2_X2 U2098 ( .A1(decode_regfile_intregs_17__13_), .A2(n13532), .ZN(n1231) );
  NAND2_X2 U2100 ( .A1(decode_regfile_intregs_17__12_), .A2(n13532), .ZN(n1232) );
  NAND2_X2 U2102 ( .A1(decode_regfile_intregs_17__11_), .A2(n13533), .ZN(n1233) );
  NAND2_X2 U2104 ( .A1(decode_regfile_intregs_17__10_), .A2(n13532), .ZN(n1234) );
  NAND2_X2 U2106 ( .A1(decode_regfile_intregs_17__0_), .A2(n13533), .ZN(n1235)
         );
  NAND2_X2 U2107 ( .A1(n1169), .A2(n800), .ZN(n1203) );
  NAND2_X2 U2109 ( .A1(decode_regfile_intregs_16__9_), .A2(n13527), .ZN(n1237)
         );
  NAND2_X2 U2111 ( .A1(decode_regfile_intregs_16__8_), .A2(n1236), .ZN(n1238)
         );
  NAND2_X2 U2113 ( .A1(decode_regfile_intregs_16__7_), .A2(n1236), .ZN(n1239)
         );
  NAND2_X2 U2115 ( .A1(decode_regfile_intregs_16__6_), .A2(n1236), .ZN(n1240)
         );
  NAND2_X2 U2117 ( .A1(decode_regfile_intregs_16__5_), .A2(n1236), .ZN(n1241)
         );
  NAND2_X2 U2119 ( .A1(decode_regfile_intregs_16__4_), .A2(n1236), .ZN(n1242)
         );
  NAND2_X2 U2121 ( .A1(decode_regfile_intregs_16__3_), .A2(n1236), .ZN(n1243)
         );
  NAND2_X2 U2123 ( .A1(decode_regfile_intregs_16__31_), .A2(n1236), .ZN(n1244)
         );
  NAND2_X2 U2125 ( .A1(decode_regfile_intregs_16__30_), .A2(n13528), .ZN(n1245) );
  NAND2_X2 U2127 ( .A1(decode_regfile_intregs_16__2_), .A2(n13528), .ZN(n1246)
         );
  NAND2_X2 U2129 ( .A1(decode_regfile_intregs_16__29_), .A2(n13528), .ZN(n1247) );
  NAND2_X2 U2131 ( .A1(decode_regfile_intregs_16__28_), .A2(n13528), .ZN(n1248) );
  NAND2_X2 U2133 ( .A1(decode_regfile_intregs_16__27_), .A2(n13528), .ZN(n1249) );
  NAND2_X2 U2135 ( .A1(decode_regfile_intregs_16__26_), .A2(n13528), .ZN(n1250) );
  NAND2_X2 U2137 ( .A1(decode_regfile_intregs_16__25_), .A2(n13528), .ZN(n1251) );
  NAND2_X2 U2139 ( .A1(decode_regfile_intregs_16__24_), .A2(n13528), .ZN(n1252) );
  NAND2_X2 U2141 ( .A1(decode_regfile_intregs_16__23_), .A2(n13528), .ZN(n1253) );
  NAND2_X2 U2143 ( .A1(decode_regfile_intregs_16__22_), .A2(n13528), .ZN(n1254) );
  NAND2_X2 U2145 ( .A1(decode_regfile_intregs_16__21_), .A2(n13528), .ZN(n1255) );
  NAND2_X2 U2147 ( .A1(decode_regfile_intregs_16__20_), .A2(n13528), .ZN(n1256) );
  NAND2_X2 U2149 ( .A1(decode_regfile_intregs_16__1_), .A2(n13528), .ZN(n1257)
         );
  NAND2_X2 U2151 ( .A1(decode_regfile_intregs_16__19_), .A2(n13528), .ZN(n1258) );
  NAND2_X2 U2153 ( .A1(decode_regfile_intregs_16__18_), .A2(n13528), .ZN(n1259) );
  NAND2_X2 U2155 ( .A1(decode_regfile_intregs_16__17_), .A2(n13528), .ZN(n1260) );
  NAND2_X2 U2157 ( .A1(decode_regfile_intregs_16__16_), .A2(n13527), .ZN(n1261) );
  NAND2_X2 U2159 ( .A1(decode_regfile_intregs_16__15_), .A2(n13527), .ZN(n1262) );
  NAND2_X2 U2161 ( .A1(decode_regfile_intregs_16__14_), .A2(n13528), .ZN(n1263) );
  NAND2_X2 U2163 ( .A1(decode_regfile_intregs_16__13_), .A2(n13527), .ZN(n1264) );
  NAND2_X2 U2165 ( .A1(decode_regfile_intregs_16__12_), .A2(n13527), .ZN(n1265) );
  NAND2_X2 U2167 ( .A1(decode_regfile_intregs_16__11_), .A2(n13528), .ZN(n1266) );
  NAND2_X2 U2169 ( .A1(decode_regfile_intregs_16__10_), .A2(n13527), .ZN(n1267) );
  NAND2_X2 U2171 ( .A1(decode_regfile_intregs_16__0_), .A2(n13528), .ZN(n1268)
         );
  NAND2_X2 U2172 ( .A1(n1169), .A2(n834), .ZN(n1236) );
  AND2_X2 U2173 ( .A1(n835), .A2(n664), .ZN(n1169) );
  NAND2_X2 U2176 ( .A1(decode_regfile_intregs_15__9_), .A2(n13522), .ZN(n1272)
         );
  NAND2_X2 U2178 ( .A1(decode_regfile_intregs_15__8_), .A2(n13524), .ZN(n1273)
         );
  NAND2_X2 U2180 ( .A1(decode_regfile_intregs_15__7_), .A2(n13524), .ZN(n1274)
         );
  NAND2_X2 U2182 ( .A1(decode_regfile_intregs_15__6_), .A2(n13524), .ZN(n1275)
         );
  NAND2_X2 U2184 ( .A1(decode_regfile_intregs_15__5_), .A2(n13524), .ZN(n1276)
         );
  NAND2_X2 U2186 ( .A1(decode_regfile_intregs_15__4_), .A2(n13524), .ZN(n1277)
         );
  NAND2_X2 U2188 ( .A1(decode_regfile_intregs_15__3_), .A2(n13524), .ZN(n1278)
         );
  NAND2_X2 U2190 ( .A1(decode_regfile_intregs_15__31_), .A2(n13524), .ZN(n1279) );
  NAND2_X2 U2192 ( .A1(decode_regfile_intregs_15__30_), .A2(n13523), .ZN(n1280) );
  NAND2_X2 U2194 ( .A1(decode_regfile_intregs_15__2_), .A2(n13523), .ZN(n1281)
         );
  NAND2_X2 U2196 ( .A1(decode_regfile_intregs_15__29_), .A2(n13523), .ZN(n1282) );
  NAND2_X2 U2198 ( .A1(decode_regfile_intregs_15__28_), .A2(n13523), .ZN(n1283) );
  NAND2_X2 U2200 ( .A1(decode_regfile_intregs_15__27_), .A2(n13523), .ZN(n1284) );
  NAND2_X2 U2202 ( .A1(decode_regfile_intregs_15__26_), .A2(n13523), .ZN(n1285) );
  NAND2_X2 U2204 ( .A1(decode_regfile_intregs_15__25_), .A2(n13523), .ZN(n1286) );
  NAND2_X2 U2206 ( .A1(decode_regfile_intregs_15__24_), .A2(n13523), .ZN(n1287) );
  NAND2_X2 U2208 ( .A1(decode_regfile_intregs_15__23_), .A2(n13523), .ZN(n1288) );
  NAND2_X2 U2210 ( .A1(decode_regfile_intregs_15__22_), .A2(n13523), .ZN(n1289) );
  NAND2_X2 U2212 ( .A1(decode_regfile_intregs_15__21_), .A2(n13523), .ZN(n1290) );
  NAND2_X2 U2214 ( .A1(decode_regfile_intregs_15__20_), .A2(n13523), .ZN(n1291) );
  NAND2_X2 U2216 ( .A1(decode_regfile_intregs_15__1_), .A2(n13523), .ZN(n1292)
         );
  NAND2_X2 U2218 ( .A1(decode_regfile_intregs_15__19_), .A2(n13523), .ZN(n1293) );
  NAND2_X2 U2220 ( .A1(decode_regfile_intregs_15__18_), .A2(n13523), .ZN(n1294) );
  NAND2_X2 U2222 ( .A1(decode_regfile_intregs_15__17_), .A2(n13523), .ZN(n1295) );
  NAND2_X2 U2224 ( .A1(decode_regfile_intregs_15__16_), .A2(n13522), .ZN(n1296) );
  NAND2_X2 U2226 ( .A1(decode_regfile_intregs_15__15_), .A2(n13522), .ZN(n1297) );
  NAND2_X2 U2228 ( .A1(decode_regfile_intregs_15__14_), .A2(n13523), .ZN(n1298) );
  NAND2_X2 U2230 ( .A1(decode_regfile_intregs_15__13_), .A2(n13522), .ZN(n1299) );
  NAND2_X2 U2232 ( .A1(decode_regfile_intregs_15__12_), .A2(n13522), .ZN(n1300) );
  NAND2_X2 U2234 ( .A1(decode_regfile_intregs_15__11_), .A2(n13523), .ZN(n1301) );
  NAND2_X2 U2236 ( .A1(decode_regfile_intregs_15__10_), .A2(n13522), .ZN(n1302) );
  NAND2_X2 U2238 ( .A1(decode_regfile_intregs_15__0_), .A2(n13523), .ZN(n1303)
         );
  NAND2_X2 U2241 ( .A1(decode_regfile_intregs_14__9_), .A2(n13517), .ZN(n1305)
         );
  NAND2_X2 U2243 ( .A1(decode_regfile_intregs_14__8_), .A2(n13519), .ZN(n1306)
         );
  NAND2_X2 U2245 ( .A1(decode_regfile_intregs_14__7_), .A2(n13519), .ZN(n1307)
         );
  NAND2_X2 U2247 ( .A1(decode_regfile_intregs_14__6_), .A2(n13519), .ZN(n1308)
         );
  NAND2_X2 U2249 ( .A1(decode_regfile_intregs_14__5_), .A2(n13519), .ZN(n1309)
         );
  NAND2_X2 U2251 ( .A1(decode_regfile_intregs_14__4_), .A2(n13519), .ZN(n1310)
         );
  NAND2_X2 U2253 ( .A1(decode_regfile_intregs_14__3_), .A2(n13519), .ZN(n1311)
         );
  NAND2_X2 U2255 ( .A1(decode_regfile_intregs_14__31_), .A2(n13519), .ZN(n1312) );
  NAND2_X2 U2257 ( .A1(decode_regfile_intregs_14__30_), .A2(n13518), .ZN(n1313) );
  NAND2_X2 U2259 ( .A1(decode_regfile_intregs_14__2_), .A2(n13518), .ZN(n1314)
         );
  NAND2_X2 U2261 ( .A1(decode_regfile_intregs_14__29_), .A2(n13518), .ZN(n1315) );
  NAND2_X2 U2263 ( .A1(decode_regfile_intregs_14__28_), .A2(n13518), .ZN(n1316) );
  NAND2_X2 U2265 ( .A1(decode_regfile_intregs_14__27_), .A2(n13518), .ZN(n1317) );
  NAND2_X2 U2267 ( .A1(decode_regfile_intregs_14__26_), .A2(n13518), .ZN(n1318) );
  NAND2_X2 U2269 ( .A1(decode_regfile_intregs_14__25_), .A2(n13518), .ZN(n1319) );
  NAND2_X2 U2271 ( .A1(decode_regfile_intregs_14__24_), .A2(n13518), .ZN(n1320) );
  NAND2_X2 U2273 ( .A1(decode_regfile_intregs_14__23_), .A2(n13518), .ZN(n1321) );
  NAND2_X2 U2275 ( .A1(decode_regfile_intregs_14__22_), .A2(n13518), .ZN(n1322) );
  NAND2_X2 U2277 ( .A1(decode_regfile_intregs_14__21_), .A2(n13518), .ZN(n1323) );
  NAND2_X2 U2279 ( .A1(decode_regfile_intregs_14__20_), .A2(n13518), .ZN(n1324) );
  NAND2_X2 U2281 ( .A1(decode_regfile_intregs_14__1_), .A2(n13518), .ZN(n1325)
         );
  NAND2_X2 U2283 ( .A1(decode_regfile_intregs_14__19_), .A2(n13518), .ZN(n1326) );
  NAND2_X2 U2285 ( .A1(decode_regfile_intregs_14__18_), .A2(n13518), .ZN(n1327) );
  NAND2_X2 U2287 ( .A1(decode_regfile_intregs_14__17_), .A2(n13518), .ZN(n1328) );
  NAND2_X2 U2289 ( .A1(decode_regfile_intregs_14__16_), .A2(n13517), .ZN(n1329) );
  NAND2_X2 U2291 ( .A1(decode_regfile_intregs_14__15_), .A2(n13517), .ZN(n1330) );
  NAND2_X2 U2293 ( .A1(decode_regfile_intregs_14__14_), .A2(n13518), .ZN(n1331) );
  NAND2_X2 U2295 ( .A1(decode_regfile_intregs_14__13_), .A2(n13517), .ZN(n1332) );
  NAND2_X2 U2297 ( .A1(decode_regfile_intregs_14__12_), .A2(n13517), .ZN(n1333) );
  NAND2_X2 U2299 ( .A1(decode_regfile_intregs_14__11_), .A2(n13518), .ZN(n1334) );
  NAND2_X2 U2301 ( .A1(decode_regfile_intregs_14__10_), .A2(n13517), .ZN(n1335) );
  NAND2_X2 U2303 ( .A1(decode_regfile_intregs_14__0_), .A2(n13518), .ZN(n1336)
         );
  NAND2_X2 U2306 ( .A1(decode_regfile_intregs_13__9_), .A2(n13512), .ZN(n1338)
         );
  NAND2_X2 U2308 ( .A1(decode_regfile_intregs_13__8_), .A2(n13514), .ZN(n1339)
         );
  NAND2_X2 U2310 ( .A1(decode_regfile_intregs_13__7_), .A2(n13514), .ZN(n1340)
         );
  NAND2_X2 U2312 ( .A1(decode_regfile_intregs_13__6_), .A2(n13514), .ZN(n1341)
         );
  NAND2_X2 U2314 ( .A1(decode_regfile_intregs_13__5_), .A2(n13514), .ZN(n1342)
         );
  NAND2_X2 U2316 ( .A1(decode_regfile_intregs_13__4_), .A2(n13514), .ZN(n1343)
         );
  NAND2_X2 U2318 ( .A1(decode_regfile_intregs_13__3_), .A2(n13514), .ZN(n1344)
         );
  NAND2_X2 U2320 ( .A1(decode_regfile_intregs_13__31_), .A2(n13514), .ZN(n1345) );
  NAND2_X2 U2322 ( .A1(decode_regfile_intregs_13__30_), .A2(n13513), .ZN(n1346) );
  NAND2_X2 U2324 ( .A1(decode_regfile_intregs_13__2_), .A2(n13513), .ZN(n1347)
         );
  NAND2_X2 U2326 ( .A1(decode_regfile_intregs_13__29_), .A2(n13513), .ZN(n1348) );
  NAND2_X2 U2328 ( .A1(decode_regfile_intregs_13__28_), .A2(n13513), .ZN(n1349) );
  NAND2_X2 U2330 ( .A1(decode_regfile_intregs_13__27_), .A2(n13513), .ZN(n1350) );
  NAND2_X2 U2332 ( .A1(decode_regfile_intregs_13__26_), .A2(n13513), .ZN(n1351) );
  NAND2_X2 U2334 ( .A1(decode_regfile_intregs_13__25_), .A2(n13513), .ZN(n1352) );
  NAND2_X2 U2336 ( .A1(decode_regfile_intregs_13__24_), .A2(n13513), .ZN(n1353) );
  NAND2_X2 U2338 ( .A1(decode_regfile_intregs_13__23_), .A2(n13513), .ZN(n1354) );
  NAND2_X2 U2340 ( .A1(decode_regfile_intregs_13__22_), .A2(n13513), .ZN(n1355) );
  NAND2_X2 U2342 ( .A1(decode_regfile_intregs_13__21_), .A2(n13513), .ZN(n1356) );
  NAND2_X2 U2344 ( .A1(decode_regfile_intregs_13__20_), .A2(n13513), .ZN(n1357) );
  NAND2_X2 U2346 ( .A1(decode_regfile_intregs_13__1_), .A2(n13513), .ZN(n1358)
         );
  NAND2_X2 U2348 ( .A1(decode_regfile_intregs_13__19_), .A2(n13513), .ZN(n1359) );
  NAND2_X2 U2350 ( .A1(decode_regfile_intregs_13__18_), .A2(n13513), .ZN(n1360) );
  NAND2_X2 U2352 ( .A1(decode_regfile_intregs_13__17_), .A2(n13513), .ZN(n1361) );
  NAND2_X2 U2354 ( .A1(decode_regfile_intregs_13__16_), .A2(n13512), .ZN(n1362) );
  NAND2_X2 U2356 ( .A1(decode_regfile_intregs_13__15_), .A2(n13512), .ZN(n1363) );
  NAND2_X2 U2358 ( .A1(decode_regfile_intregs_13__14_), .A2(n13513), .ZN(n1364) );
  NAND2_X2 U2360 ( .A1(decode_regfile_intregs_13__13_), .A2(n13512), .ZN(n1365) );
  NAND2_X2 U2362 ( .A1(decode_regfile_intregs_13__12_), .A2(n13512), .ZN(n1366) );
  NAND2_X2 U2364 ( .A1(decode_regfile_intregs_13__11_), .A2(n13513), .ZN(n1367) );
  NAND2_X2 U2366 ( .A1(decode_regfile_intregs_13__10_), .A2(n13512), .ZN(n1368) );
  NAND2_X2 U2368 ( .A1(decode_regfile_intregs_13__0_), .A2(n13513), .ZN(n1369)
         );
  AND2_X2 U2370 ( .A1(n1370), .A2(n800), .ZN(n460) );
  NAND2_X2 U2372 ( .A1(decode_regfile_intregs_12__9_), .A2(n13507), .ZN(n1372)
         );
  NAND2_X2 U2374 ( .A1(decode_regfile_intregs_12__8_), .A2(n13509), .ZN(n1373)
         );
  NAND2_X2 U2376 ( .A1(decode_regfile_intregs_12__7_), .A2(n13509), .ZN(n1374)
         );
  NAND2_X2 U2378 ( .A1(decode_regfile_intregs_12__6_), .A2(n13509), .ZN(n1375)
         );
  NAND2_X2 U2380 ( .A1(decode_regfile_intregs_12__5_), .A2(n13509), .ZN(n1376)
         );
  NAND2_X2 U2382 ( .A1(decode_regfile_intregs_12__4_), .A2(n13509), .ZN(n1377)
         );
  NAND2_X2 U2384 ( .A1(decode_regfile_intregs_12__3_), .A2(n13509), .ZN(n1378)
         );
  NAND2_X2 U2386 ( .A1(decode_regfile_intregs_12__31_), .A2(n13509), .ZN(n1379) );
  NAND2_X2 U2388 ( .A1(decode_regfile_intregs_12__30_), .A2(n13508), .ZN(n1380) );
  NAND2_X2 U2390 ( .A1(decode_regfile_intregs_12__2_), .A2(n13508), .ZN(n1381)
         );
  NAND2_X2 U2392 ( .A1(decode_regfile_intregs_12__29_), .A2(n13508), .ZN(n1382) );
  NAND2_X2 U2394 ( .A1(decode_regfile_intregs_12__28_), .A2(n13508), .ZN(n1383) );
  NAND2_X2 U2396 ( .A1(decode_regfile_intregs_12__27_), .A2(n13508), .ZN(n1384) );
  NAND2_X2 U2398 ( .A1(decode_regfile_intregs_12__26_), .A2(n13508), .ZN(n1385) );
  NAND2_X2 U2400 ( .A1(decode_regfile_intregs_12__25_), .A2(n13508), .ZN(n1386) );
  NAND2_X2 U2402 ( .A1(decode_regfile_intregs_12__24_), .A2(n13508), .ZN(n1387) );
  NAND2_X2 U2404 ( .A1(decode_regfile_intregs_12__23_), .A2(n13508), .ZN(n1388) );
  NAND2_X2 U2406 ( .A1(decode_regfile_intregs_12__22_), .A2(n13508), .ZN(n1389) );
  NAND2_X2 U2408 ( .A1(decode_regfile_intregs_12__21_), .A2(n13508), .ZN(n1390) );
  NAND2_X2 U2410 ( .A1(decode_regfile_intregs_12__20_), .A2(n13508), .ZN(n1391) );
  NAND2_X2 U2412 ( .A1(decode_regfile_intregs_12__1_), .A2(n13508), .ZN(n1392)
         );
  NAND2_X2 U2414 ( .A1(decode_regfile_intregs_12__19_), .A2(n13508), .ZN(n1393) );
  NAND2_X2 U2416 ( .A1(decode_regfile_intregs_12__18_), .A2(n13508), .ZN(n1394) );
  NAND2_X2 U2418 ( .A1(decode_regfile_intregs_12__17_), .A2(n13508), .ZN(n1395) );
  NAND2_X2 U2420 ( .A1(decode_regfile_intregs_12__16_), .A2(n13507), .ZN(n1396) );
  NAND2_X2 U2422 ( .A1(decode_regfile_intregs_12__15_), .A2(n13507), .ZN(n1397) );
  NAND2_X2 U2424 ( .A1(decode_regfile_intregs_12__14_), .A2(n13508), .ZN(n1398) );
  NAND2_X2 U2426 ( .A1(decode_regfile_intregs_12__13_), .A2(n13507), .ZN(n1399) );
  NAND2_X2 U2428 ( .A1(decode_regfile_intregs_12__12_), .A2(n13507), .ZN(n1400) );
  NAND2_X2 U2430 ( .A1(decode_regfile_intregs_12__11_), .A2(n13508), .ZN(n1401) );
  NAND2_X2 U2432 ( .A1(decode_regfile_intregs_12__10_), .A2(n13507), .ZN(n1402) );
  NAND2_X2 U2434 ( .A1(decode_regfile_intregs_12__0_), .A2(n13508), .ZN(n1403)
         );
  NAND2_X2 U2437 ( .A1(decode_regfile_intregs_11__9_), .A2(n13502), .ZN(n1405)
         );
  NAND2_X2 U2439 ( .A1(decode_regfile_intregs_11__8_), .A2(n13504), .ZN(n1406)
         );
  NAND2_X2 U2441 ( .A1(decode_regfile_intregs_11__7_), .A2(n13504), .ZN(n1407)
         );
  NAND2_X2 U2443 ( .A1(decode_regfile_intregs_11__6_), .A2(n13504), .ZN(n1408)
         );
  NAND2_X2 U2445 ( .A1(decode_regfile_intregs_11__5_), .A2(n13504), .ZN(n1409)
         );
  NAND2_X2 U2447 ( .A1(decode_regfile_intregs_11__4_), .A2(n13504), .ZN(n1410)
         );
  NAND2_X2 U2449 ( .A1(decode_regfile_intregs_11__3_), .A2(n13504), .ZN(n1411)
         );
  NAND2_X2 U2451 ( .A1(decode_regfile_intregs_11__31_), .A2(n13504), .ZN(n1412) );
  NAND2_X2 U2453 ( .A1(decode_regfile_intregs_11__30_), .A2(n13503), .ZN(n1413) );
  NAND2_X2 U2455 ( .A1(decode_regfile_intregs_11__2_), .A2(n13503), .ZN(n1414)
         );
  NAND2_X2 U2457 ( .A1(decode_regfile_intregs_11__29_), .A2(n13503), .ZN(n1415) );
  NAND2_X2 U2459 ( .A1(decode_regfile_intregs_11__28_), .A2(n13503), .ZN(n1416) );
  NAND2_X2 U2461 ( .A1(decode_regfile_intregs_11__27_), .A2(n13503), .ZN(n1417) );
  NAND2_X2 U2463 ( .A1(decode_regfile_intregs_11__26_), .A2(n13503), .ZN(n1418) );
  NAND2_X2 U2465 ( .A1(decode_regfile_intregs_11__25_), .A2(n13503), .ZN(n1419) );
  NAND2_X2 U2467 ( .A1(decode_regfile_intregs_11__24_), .A2(n13503), .ZN(n1420) );
  NAND2_X2 U2469 ( .A1(decode_regfile_intregs_11__23_), .A2(n13503), .ZN(n1421) );
  NAND2_X2 U2471 ( .A1(decode_regfile_intregs_11__22_), .A2(n13503), .ZN(n1422) );
  NAND2_X2 U2473 ( .A1(decode_regfile_intregs_11__21_), .A2(n13503), .ZN(n1423) );
  NAND2_X2 U2475 ( .A1(decode_regfile_intregs_11__20_), .A2(n13503), .ZN(n1424) );
  NAND2_X2 U2477 ( .A1(decode_regfile_intregs_11__1_), .A2(n13503), .ZN(n1425)
         );
  NAND2_X2 U2479 ( .A1(decode_regfile_intregs_11__19_), .A2(n13503), .ZN(n1426) );
  NAND2_X2 U2481 ( .A1(decode_regfile_intregs_11__18_), .A2(n13503), .ZN(n1427) );
  NAND2_X2 U2483 ( .A1(decode_regfile_intregs_11__17_), .A2(n13503), .ZN(n1428) );
  NAND2_X2 U2485 ( .A1(decode_regfile_intregs_11__16_), .A2(n13502), .ZN(n1429) );
  NAND2_X2 U2487 ( .A1(decode_regfile_intregs_11__15_), .A2(n13502), .ZN(n1430) );
  NAND2_X2 U2489 ( .A1(decode_regfile_intregs_11__14_), .A2(n13503), .ZN(n1431) );
  NAND2_X2 U2491 ( .A1(decode_regfile_intregs_11__13_), .A2(n13502), .ZN(n1432) );
  NAND2_X2 U2493 ( .A1(decode_regfile_intregs_11__12_), .A2(n13502), .ZN(n1433) );
  NAND2_X2 U2495 ( .A1(decode_regfile_intregs_11__11_), .A2(n13503), .ZN(n1434) );
  NAND2_X2 U2497 ( .A1(decode_regfile_intregs_11__10_), .A2(n13502), .ZN(n1435) );
  NAND2_X2 U2499 ( .A1(decode_regfile_intregs_11__0_), .A2(n13503), .ZN(n1436)
         );
  AND2_X2 U2501 ( .A1(n699), .A2(n1370), .ZN(n529) );
  NAND2_X2 U2503 ( .A1(decode_regfile_intregs_10__9_), .A2(n13497), .ZN(n1438)
         );
  NAND2_X2 U2505 ( .A1(decode_regfile_intregs_10__8_), .A2(n13499), .ZN(n1439)
         );
  NAND2_X2 U2507 ( .A1(decode_regfile_intregs_10__7_), .A2(n13499), .ZN(n1440)
         );
  NAND2_X2 U2509 ( .A1(decode_regfile_intregs_10__6_), .A2(n13499), .ZN(n1441)
         );
  NAND2_X2 U2511 ( .A1(decode_regfile_intregs_10__5_), .A2(n13499), .ZN(n1442)
         );
  NAND2_X2 U2513 ( .A1(decode_regfile_intregs_10__4_), .A2(n13499), .ZN(n1443)
         );
  NAND2_X2 U2515 ( .A1(decode_regfile_intregs_10__3_), .A2(n13499), .ZN(n1444)
         );
  NAND2_X2 U2517 ( .A1(decode_regfile_intregs_10__31_), .A2(n13499), .ZN(n1445) );
  NAND2_X2 U2519 ( .A1(decode_regfile_intregs_10__30_), .A2(n13498), .ZN(n1446) );
  NAND2_X2 U2521 ( .A1(decode_regfile_intregs_10__2_), .A2(n13498), .ZN(n1447)
         );
  NAND2_X2 U2523 ( .A1(decode_regfile_intregs_10__29_), .A2(n13498), .ZN(n1448) );
  NAND2_X2 U2525 ( .A1(decode_regfile_intregs_10__28_), .A2(n13498), .ZN(n1449) );
  NAND2_X2 U2527 ( .A1(decode_regfile_intregs_10__27_), .A2(n13498), .ZN(n1450) );
  NAND2_X2 U2529 ( .A1(decode_regfile_intregs_10__26_), .A2(n13498), .ZN(n1451) );
  NAND2_X2 U2531 ( .A1(decode_regfile_intregs_10__25_), .A2(n13498), .ZN(n1452) );
  NAND2_X2 U2533 ( .A1(decode_regfile_intregs_10__24_), .A2(n13498), .ZN(n1453) );
  NAND2_X2 U2535 ( .A1(decode_regfile_intregs_10__23_), .A2(n13498), .ZN(n1454) );
  NAND2_X2 U2537 ( .A1(decode_regfile_intregs_10__22_), .A2(n13498), .ZN(n1455) );
  NAND2_X2 U2539 ( .A1(decode_regfile_intregs_10__21_), .A2(n13498), .ZN(n1456) );
  NAND2_X2 U2541 ( .A1(decode_regfile_intregs_10__20_), .A2(n13498), .ZN(n1457) );
  NAND2_X2 U2543 ( .A1(decode_regfile_intregs_10__1_), .A2(n13498), .ZN(n1458)
         );
  NAND2_X2 U2545 ( .A1(decode_regfile_intregs_10__19_), .A2(n13498), .ZN(n1459) );
  NAND2_X2 U2547 ( .A1(decode_regfile_intregs_10__18_), .A2(n13498), .ZN(n1460) );
  NAND2_X2 U2549 ( .A1(decode_regfile_intregs_10__17_), .A2(n13498), .ZN(n1461) );
  NAND2_X2 U2551 ( .A1(decode_regfile_intregs_10__16_), .A2(n13497), .ZN(n1462) );
  NAND2_X2 U2553 ( .A1(decode_regfile_intregs_10__15_), .A2(n13497), .ZN(n1463) );
  NAND2_X2 U2555 ( .A1(decode_regfile_intregs_10__14_), .A2(n13498), .ZN(n1464) );
  NAND2_X2 U2557 ( .A1(decode_regfile_intregs_10__13_), .A2(n13497), .ZN(n1465) );
  NAND2_X2 U2559 ( .A1(decode_regfile_intregs_10__12_), .A2(n13497), .ZN(n1466) );
  NAND2_X2 U2561 ( .A1(decode_regfile_intregs_10__11_), .A2(n13498), .ZN(n1467) );
  NAND2_X2 U2563 ( .A1(decode_regfile_intregs_10__10_), .A2(n13497), .ZN(n1468) );
  NAND2_X2 U2565 ( .A1(decode_regfile_intregs_10__0_), .A2(n13498), .ZN(n1469)
         );
  AND2_X2 U2567 ( .A1(n733), .A2(n1370), .ZN(n564) );
  NAND2_X2 U2569 ( .A1(decode_regfile_intregs_0__9_), .A2(n13492), .ZN(n1471)
         );
  AOI22_X2 U2570 ( .A1(decode_regfile_N154), .A2(n13489), .B1(n16552), .B2(
        n13487), .ZN(n395) );
  NAND2_X2 U2572 ( .A1(decode_regfile_intregs_0__8_), .A2(n13494), .ZN(n1474)
         );
  AOI22_X2 U2573 ( .A1(decode_regfile_N155), .A2(n13488), .B1(n16553), .B2(
        n13486), .ZN(n398) );
  NAND2_X2 U2575 ( .A1(decode_regfile_intregs_0__7_), .A2(n13494), .ZN(n1475)
         );
  AOI22_X2 U2576 ( .A1(decode_regfile_N156), .A2(n13488), .B1(n16554), .B2(
        n13486), .ZN(n400) );
  NAND2_X2 U2578 ( .A1(decode_regfile_intregs_0__6_), .A2(n13494), .ZN(n1476)
         );
  AOI22_X2 U2579 ( .A1(decode_regfile_N157), .A2(n13488), .B1(n16555), .B2(
        n13486), .ZN(n402) );
  NAND2_X2 U2581 ( .A1(decode_regfile_intregs_0__5_), .A2(n13494), .ZN(n1477)
         );
  AOI22_X2 U2582 ( .A1(decode_regfile_N158), .A2(n13488), .B1(n16556), .B2(
        n13486), .ZN(n404) );
  NAND2_X2 U2584 ( .A1(decode_regfile_intregs_0__4_), .A2(n13494), .ZN(n1478)
         );
  AOI22_X2 U2585 ( .A1(decode_regfile_N159), .A2(n13488), .B1(n16557), .B2(
        n13486), .ZN(n406) );
  NAND2_X2 U2587 ( .A1(decode_regfile_intregs_0__3_), .A2(n13494), .ZN(n1479)
         );
  AOI22_X2 U2588 ( .A1(decode_regfile_N160), .A2(n13488), .B1(n16558), .B2(
        n13486), .ZN(n408) );
  NAND2_X2 U2590 ( .A1(decode_regfile_intregs_0__31_), .A2(n13494), .ZN(n1480)
         );
  AOI22_X2 U2591 ( .A1(decode_regfile_N132), .A2(n13488), .B1(n16559), .B2(
        n13486), .ZN(n410) );
  NAND2_X2 U2593 ( .A1(decode_regfile_intregs_0__30_), .A2(n13493), .ZN(n1481)
         );
  AOI22_X2 U2594 ( .A1(decode_regfile_N133), .A2(n13488), .B1(n16560), .B2(
        n13486), .ZN(n412) );
  NAND2_X2 U2596 ( .A1(decode_regfile_intregs_0__2_), .A2(n13493), .ZN(n1482)
         );
  AOI22_X2 U2597 ( .A1(decode_regfile_N161), .A2(n13488), .B1(n16561), .B2(
        n13486), .ZN(n414) );
  NAND2_X2 U2599 ( .A1(decode_regfile_intregs_0__29_), .A2(n13493), .ZN(n1483)
         );
  AOI22_X2 U2600 ( .A1(decode_regfile_N134), .A2(n13488), .B1(n16562), .B2(
        n13486), .ZN(n416) );
  NAND2_X2 U2602 ( .A1(decode_regfile_intregs_0__28_), .A2(n13493), .ZN(n1484)
         );
  AOI22_X2 U2603 ( .A1(decode_regfile_N135), .A2(n13488), .B1(n16563), .B2(
        n13486), .ZN(n418) );
  NAND2_X2 U2605 ( .A1(decode_regfile_intregs_0__27_), .A2(n13493), .ZN(n1485)
         );
  AOI22_X2 U2606 ( .A1(decode_regfile_N136), .A2(n13488), .B1(n16564), .B2(
        n13486), .ZN(n420) );
  NAND2_X2 U2608 ( .A1(decode_regfile_intregs_0__26_), .A2(n13493), .ZN(n1486)
         );
  AOI22_X2 U2609 ( .A1(decode_regfile_N137), .A2(n13488), .B1(n16565), .B2(
        n13486), .ZN(n422) );
  NAND2_X2 U2611 ( .A1(decode_regfile_intregs_0__25_), .A2(n13493), .ZN(n1487)
         );
  AOI22_X2 U2612 ( .A1(decode_regfile_N138), .A2(n13488), .B1(n16566), .B2(
        n13486), .ZN(n424) );
  NAND2_X2 U2614 ( .A1(decode_regfile_intregs_0__24_), .A2(n13493), .ZN(n1488)
         );
  AOI22_X2 U2615 ( .A1(decode_regfile_N139), .A2(n13488), .B1(n16567), .B2(
        n13486), .ZN(n426) );
  NAND2_X2 U2617 ( .A1(decode_regfile_intregs_0__23_), .A2(n13493), .ZN(n1489)
         );
  AOI22_X2 U2618 ( .A1(decode_regfile_N140), .A2(n13489), .B1(n16568), .B2(
        n13487), .ZN(n428) );
  NAND2_X2 U2620 ( .A1(decode_regfile_intregs_0__22_), .A2(n13493), .ZN(n1490)
         );
  AOI22_X2 U2621 ( .A1(decode_regfile_N141), .A2(n13489), .B1(n16569), .B2(
        n13487), .ZN(n430) );
  NAND2_X2 U2623 ( .A1(decode_regfile_intregs_0__21_), .A2(n13493), .ZN(n1491)
         );
  AOI22_X2 U2624 ( .A1(decode_regfile_N142), .A2(n13489), .B1(n16570), .B2(
        n13487), .ZN(n432) );
  NAND2_X2 U2626 ( .A1(decode_regfile_intregs_0__20_), .A2(n13493), .ZN(n1492)
         );
  AOI22_X2 U2627 ( .A1(decode_regfile_N143), .A2(n13489), .B1(n16571), .B2(
        n13487), .ZN(n434) );
  NAND2_X2 U2629 ( .A1(decode_regfile_intregs_0__1_), .A2(n13493), .ZN(n1493)
         );
  AOI22_X2 U2630 ( .A1(decode_regfile_N162), .A2(n13489), .B1(n16572), .B2(
        n13487), .ZN(n436) );
  NAND2_X2 U2632 ( .A1(decode_regfile_intregs_0__19_), .A2(n13493), .ZN(n1494)
         );
  AOI22_X2 U2633 ( .A1(decode_regfile_N144), .A2(n13489), .B1(n16255), .B2(
        n13487), .ZN(n438) );
  NAND2_X2 U2635 ( .A1(decode_regfile_intregs_0__18_), .A2(n13493), .ZN(n1495)
         );
  AOI22_X2 U2636 ( .A1(decode_regfile_N145), .A2(n13489), .B1(n16573), .B2(
        n13487), .ZN(n440) );
  NAND2_X2 U2638 ( .A1(decode_regfile_intregs_0__17_), .A2(n13493), .ZN(n1496)
         );
  AOI22_X2 U2639 ( .A1(decode_regfile_N146), .A2(n13489), .B1(n16574), .B2(
        n13487), .ZN(n442) );
  NAND2_X2 U2641 ( .A1(decode_regfile_intregs_0__16_), .A2(n13492), .ZN(n1497)
         );
  AOI22_X2 U2642 ( .A1(decode_regfile_N147), .A2(n13489), .B1(n16575), .B2(
        n13487), .ZN(n444) );
  NAND2_X2 U2644 ( .A1(decode_regfile_intregs_0__15_), .A2(n13492), .ZN(n1498)
         );
  AOI22_X2 U2645 ( .A1(decode_regfile_N148), .A2(n13489), .B1(n16576), .B2(
        n13487), .ZN(n446) );
  NAND2_X2 U2647 ( .A1(decode_regfile_intregs_0__14_), .A2(n13493), .ZN(n1499)
         );
  AOI22_X2 U2648 ( .A1(decode_regfile_N149), .A2(n13489), .B1(n16577), .B2(
        n13487), .ZN(n448) );
  NAND2_X2 U2650 ( .A1(decode_regfile_intregs_0__13_), .A2(n13492), .ZN(n1500)
         );
  AOI22_X2 U2651 ( .A1(decode_regfile_N150), .A2(n13489), .B1(n16578), .B2(
        n13487), .ZN(n450) );
  NAND2_X2 U2653 ( .A1(decode_regfile_intregs_0__12_), .A2(n13492), .ZN(n1501)
         );
  AOI22_X2 U2654 ( .A1(decode_regfile_N151), .A2(n13489), .B1(n16579), .B2(
        n13487), .ZN(n452) );
  NAND2_X2 U2656 ( .A1(decode_regfile_intregs_0__11_), .A2(n13493), .ZN(n1502)
         );
  AOI22_X2 U2657 ( .A1(decode_regfile_N152), .A2(n13489), .B1(n16580), .B2(
        n13487), .ZN(n454) );
  NAND2_X2 U2659 ( .A1(decode_regfile_intregs_0__10_), .A2(n13492), .ZN(n1503)
         );
  AOI22_X2 U2660 ( .A1(decode_regfile_N153), .A2(n13489), .B1(n16581), .B2(
        n13487), .ZN(n456) );
  NAND2_X2 U2662 ( .A1(decode_regfile_intregs_0__0_), .A2(n13493), .ZN(n1504)
         );
  AND2_X2 U2664 ( .A1(n834), .A2(n1370), .ZN(n495) );
  AOI22_X2 U2667 ( .A1(decode_regfile_N163), .A2(n13488), .B1(n16582), .B2(
        n13486), .ZN(n458) );
  NAND2_X2 U2671 ( .A1(decode_regfile_fpregs_9__9_), .A2(n13480), .ZN(n1508)
         );
  NAND2_X2 U2673 ( .A1(decode_regfile_fpregs_9__8_), .A2(n1507), .ZN(n1510) );
  NAND2_X2 U2675 ( .A1(decode_regfile_fpregs_9__7_), .A2(n1507), .ZN(n1512) );
  NAND2_X2 U2677 ( .A1(decode_regfile_fpregs_9__6_), .A2(n1507), .ZN(n1514) );
  NAND2_X2 U2679 ( .A1(decode_regfile_fpregs_9__5_), .A2(n1507), .ZN(n1516) );
  NAND2_X2 U2681 ( .A1(decode_regfile_fpregs_9__4_), .A2(n1507), .ZN(n1518) );
  NAND2_X2 U2683 ( .A1(decode_regfile_fpregs_9__3_), .A2(n1507), .ZN(n1520) );
  NAND2_X2 U2685 ( .A1(decode_regfile_fpregs_9__31_), .A2(n1507), .ZN(n1522)
         );
  NAND2_X2 U2687 ( .A1(decode_regfile_fpregs_9__30_), .A2(n13481), .ZN(n1524)
         );
  NAND2_X2 U2689 ( .A1(decode_regfile_fpregs_9__2_), .A2(n13481), .ZN(n1526)
         );
  NAND2_X2 U2691 ( .A1(decode_regfile_fpregs_9__29_), .A2(n13481), .ZN(n1528)
         );
  NAND2_X2 U2693 ( .A1(decode_regfile_fpregs_9__28_), .A2(n13481), .ZN(n1530)
         );
  NAND2_X2 U2695 ( .A1(decode_regfile_fpregs_9__27_), .A2(n13481), .ZN(n1532)
         );
  NAND2_X2 U2697 ( .A1(decode_regfile_fpregs_9__26_), .A2(n13481), .ZN(n1534)
         );
  NAND2_X2 U2699 ( .A1(decode_regfile_fpregs_9__25_), .A2(n13481), .ZN(n1536)
         );
  NAND2_X2 U2701 ( .A1(decode_regfile_fpregs_9__24_), .A2(n13481), .ZN(n1538)
         );
  NAND2_X2 U2703 ( .A1(decode_regfile_fpregs_9__23_), .A2(n13481), .ZN(n1540)
         );
  NAND2_X2 U2705 ( .A1(decode_regfile_fpregs_9__22_), .A2(n13481), .ZN(n1542)
         );
  NAND2_X2 U2707 ( .A1(decode_regfile_fpregs_9__21_), .A2(n13481), .ZN(n1544)
         );
  NAND2_X2 U2709 ( .A1(decode_regfile_fpregs_9__20_), .A2(n13481), .ZN(n1546)
         );
  NAND2_X2 U2711 ( .A1(decode_regfile_fpregs_9__1_), .A2(n13481), .ZN(n1548)
         );
  NAND2_X2 U2713 ( .A1(decode_regfile_fpregs_9__19_), .A2(n13481), .ZN(n1550)
         );
  NAND2_X2 U2715 ( .A1(decode_regfile_fpregs_9__18_), .A2(n13481), .ZN(n1552)
         );
  NAND2_X2 U2717 ( .A1(decode_regfile_fpregs_9__17_), .A2(n13481), .ZN(n1554)
         );
  NAND2_X2 U2719 ( .A1(decode_regfile_fpregs_9__16_), .A2(n13480), .ZN(n1556)
         );
  NAND2_X2 U2721 ( .A1(decode_regfile_fpregs_9__15_), .A2(n13480), .ZN(n1558)
         );
  NAND2_X2 U2723 ( .A1(decode_regfile_fpregs_9__14_), .A2(n13481), .ZN(n1560)
         );
  NAND2_X2 U2725 ( .A1(decode_regfile_fpregs_9__13_), .A2(n13480), .ZN(n1562)
         );
  NAND2_X2 U2727 ( .A1(decode_regfile_fpregs_9__12_), .A2(n13480), .ZN(n1564)
         );
  NAND2_X2 U2729 ( .A1(decode_regfile_fpregs_9__11_), .A2(n13481), .ZN(n1566)
         );
  NAND2_X2 U2731 ( .A1(decode_regfile_fpregs_9__10_), .A2(n13480), .ZN(n1568)
         );
  NAND2_X2 U2733 ( .A1(decode_regfile_fpregs_9__0_), .A2(n13481), .ZN(n1570)
         );
  NAND2_X2 U2734 ( .A1(n1571), .A2(n800), .ZN(n1507) );
  NAND2_X2 U2736 ( .A1(decode_regfile_fpregs_8__9_), .A2(n13382), .ZN(n1573)
         );
  NAND2_X2 U2738 ( .A1(decode_regfile_fpregs_8__8_), .A2(n1572), .ZN(n1574) );
  NAND2_X2 U2740 ( .A1(decode_regfile_fpregs_8__7_), .A2(n1572), .ZN(n1575) );
  NAND2_X2 U2742 ( .A1(decode_regfile_fpregs_8__6_), .A2(n1572), .ZN(n1576) );
  NAND2_X2 U2744 ( .A1(decode_regfile_fpregs_8__5_), .A2(n1572), .ZN(n1577) );
  NAND2_X2 U2746 ( .A1(decode_regfile_fpregs_8__4_), .A2(n1572), .ZN(n1578) );
  NAND2_X2 U2748 ( .A1(decode_regfile_fpregs_8__3_), .A2(n1572), .ZN(n1579) );
  NAND2_X2 U2750 ( .A1(decode_regfile_fpregs_8__31_), .A2(n1572), .ZN(n1580)
         );
  NAND2_X2 U2752 ( .A1(decode_regfile_fpregs_8__30_), .A2(n13383), .ZN(n1581)
         );
  NAND2_X2 U2754 ( .A1(decode_regfile_fpregs_8__2_), .A2(n13383), .ZN(n1582)
         );
  NAND2_X2 U2756 ( .A1(decode_regfile_fpregs_8__29_), .A2(n13383), .ZN(n1583)
         );
  NAND2_X2 U2758 ( .A1(decode_regfile_fpregs_8__28_), .A2(n13383), .ZN(n1584)
         );
  NAND2_X2 U2760 ( .A1(decode_regfile_fpregs_8__27_), .A2(n13383), .ZN(n1585)
         );
  NAND2_X2 U2762 ( .A1(decode_regfile_fpregs_8__26_), .A2(n13383), .ZN(n1586)
         );
  NAND2_X2 U2764 ( .A1(decode_regfile_fpregs_8__25_), .A2(n13383), .ZN(n1587)
         );
  NAND2_X2 U2766 ( .A1(decode_regfile_fpregs_8__24_), .A2(n13383), .ZN(n1588)
         );
  NAND2_X2 U2768 ( .A1(decode_regfile_fpregs_8__23_), .A2(n13383), .ZN(n1589)
         );
  NAND2_X2 U2770 ( .A1(decode_regfile_fpregs_8__22_), .A2(n13383), .ZN(n1590)
         );
  NAND2_X2 U2772 ( .A1(decode_regfile_fpregs_8__21_), .A2(n13383), .ZN(n1591)
         );
  NAND2_X2 U2774 ( .A1(decode_regfile_fpregs_8__20_), .A2(n13383), .ZN(n1592)
         );
  NAND2_X2 U2776 ( .A1(decode_regfile_fpregs_8__1_), .A2(n13383), .ZN(n1593)
         );
  NAND2_X2 U2778 ( .A1(decode_regfile_fpregs_8__19_), .A2(n13383), .ZN(n1594)
         );
  NAND2_X2 U2780 ( .A1(decode_regfile_fpregs_8__18_), .A2(n13383), .ZN(n1595)
         );
  NAND2_X2 U2782 ( .A1(decode_regfile_fpregs_8__17_), .A2(n13383), .ZN(n1596)
         );
  NAND2_X2 U2784 ( .A1(decode_regfile_fpregs_8__16_), .A2(n13382), .ZN(n1597)
         );
  NAND2_X2 U2786 ( .A1(decode_regfile_fpregs_8__15_), .A2(n13382), .ZN(n1598)
         );
  NAND2_X2 U2788 ( .A1(decode_regfile_fpregs_8__14_), .A2(n13383), .ZN(n1599)
         );
  NAND2_X2 U2790 ( .A1(decode_regfile_fpregs_8__13_), .A2(n13382), .ZN(n1600)
         );
  NAND2_X2 U2792 ( .A1(decode_regfile_fpregs_8__12_), .A2(n13382), .ZN(n1601)
         );
  NAND2_X2 U2794 ( .A1(decode_regfile_fpregs_8__11_), .A2(n13383), .ZN(n1602)
         );
  NAND2_X2 U2796 ( .A1(decode_regfile_fpregs_8__10_), .A2(n13382), .ZN(n1603)
         );
  NAND2_X2 U2798 ( .A1(decode_regfile_fpregs_8__0_), .A2(n13383), .ZN(n1604)
         );
  NAND2_X2 U2799 ( .A1(n1571), .A2(n834), .ZN(n1572) );
  NAND2_X2 U2801 ( .A1(decode_regfile_fpregs_7__9_), .A2(n13377), .ZN(n1606)
         );
  NAND2_X2 U2803 ( .A1(decode_regfile_fpregs_7__8_), .A2(n13379), .ZN(n1607)
         );
  NAND2_X2 U2805 ( .A1(decode_regfile_fpregs_7__7_), .A2(n13379), .ZN(n1608)
         );
  NAND2_X2 U2807 ( .A1(decode_regfile_fpregs_7__6_), .A2(n13379), .ZN(n1609)
         );
  NAND2_X2 U2809 ( .A1(decode_regfile_fpregs_7__5_), .A2(n13379), .ZN(n1610)
         );
  NAND2_X2 U2811 ( .A1(decode_regfile_fpregs_7__4_), .A2(n13379), .ZN(n1611)
         );
  NAND2_X2 U2813 ( .A1(decode_regfile_fpregs_7__3_), .A2(n13379), .ZN(n1612)
         );
  NAND2_X2 U2815 ( .A1(decode_regfile_fpregs_7__31_), .A2(n13379), .ZN(n1613)
         );
  NAND2_X2 U2817 ( .A1(decode_regfile_fpregs_7__30_), .A2(n13378), .ZN(n1614)
         );
  NAND2_X2 U2819 ( .A1(decode_regfile_fpregs_7__2_), .A2(n13378), .ZN(n1615)
         );
  NAND2_X2 U2821 ( .A1(decode_regfile_fpregs_7__29_), .A2(n13378), .ZN(n1616)
         );
  NAND2_X2 U2823 ( .A1(decode_regfile_fpregs_7__28_), .A2(n13378), .ZN(n1617)
         );
  NAND2_X2 U2825 ( .A1(decode_regfile_fpregs_7__27_), .A2(n13378), .ZN(n1618)
         );
  NAND2_X2 U2827 ( .A1(decode_regfile_fpregs_7__26_), .A2(n13378), .ZN(n1619)
         );
  NAND2_X2 U2829 ( .A1(decode_regfile_fpregs_7__25_), .A2(n13378), .ZN(n1620)
         );
  NAND2_X2 U2831 ( .A1(decode_regfile_fpregs_7__24_), .A2(n13378), .ZN(n1621)
         );
  NAND2_X2 U2833 ( .A1(decode_regfile_fpregs_7__23_), .A2(n13378), .ZN(n1622)
         );
  NAND2_X2 U2835 ( .A1(decode_regfile_fpregs_7__22_), .A2(n13378), .ZN(n1623)
         );
  NAND2_X2 U2837 ( .A1(decode_regfile_fpregs_7__21_), .A2(n13378), .ZN(n1624)
         );
  NAND2_X2 U2839 ( .A1(decode_regfile_fpregs_7__20_), .A2(n13378), .ZN(n1625)
         );
  NAND2_X2 U2841 ( .A1(decode_regfile_fpregs_7__1_), .A2(n13378), .ZN(n1626)
         );
  NAND2_X2 U2843 ( .A1(decode_regfile_fpregs_7__19_), .A2(n13378), .ZN(n1627)
         );
  NAND2_X2 U2845 ( .A1(decode_regfile_fpregs_7__18_), .A2(n13378), .ZN(n1628)
         );
  NAND2_X2 U2847 ( .A1(decode_regfile_fpregs_7__17_), .A2(n13378), .ZN(n1629)
         );
  NAND2_X2 U2849 ( .A1(decode_regfile_fpregs_7__16_), .A2(n13377), .ZN(n1630)
         );
  NAND2_X2 U2851 ( .A1(decode_regfile_fpregs_7__15_), .A2(n13377), .ZN(n1631)
         );
  NAND2_X2 U2853 ( .A1(decode_regfile_fpregs_7__14_), .A2(n13378), .ZN(n1632)
         );
  NAND2_X2 U2855 ( .A1(decode_regfile_fpregs_7__13_), .A2(n13377), .ZN(n1633)
         );
  NAND2_X2 U2857 ( .A1(decode_regfile_fpregs_7__12_), .A2(n13377), .ZN(n1634)
         );
  NAND2_X2 U2859 ( .A1(decode_regfile_fpregs_7__11_), .A2(n13378), .ZN(n1635)
         );
  NAND2_X2 U2861 ( .A1(decode_regfile_fpregs_7__10_), .A2(n13377), .ZN(n1636)
         );
  NAND2_X2 U2863 ( .A1(decode_regfile_fpregs_7__0_), .A2(n13378), .ZN(n1637)
         );
  NAND2_X2 U2866 ( .A1(decode_regfile_fpregs_6__9_), .A2(n13372), .ZN(n1640)
         );
  NAND2_X2 U2868 ( .A1(decode_regfile_fpregs_6__8_), .A2(n13374), .ZN(n1641)
         );
  NAND2_X2 U2870 ( .A1(decode_regfile_fpregs_6__7_), .A2(n13374), .ZN(n1642)
         );
  NAND2_X2 U2872 ( .A1(decode_regfile_fpregs_6__6_), .A2(n13374), .ZN(n1643)
         );
  NAND2_X2 U2874 ( .A1(decode_regfile_fpregs_6__5_), .A2(n13374), .ZN(n1644)
         );
  NAND2_X2 U2876 ( .A1(decode_regfile_fpregs_6__4_), .A2(n13374), .ZN(n1645)
         );
  NAND2_X2 U2878 ( .A1(decode_regfile_fpregs_6__3_), .A2(n13374), .ZN(n1646)
         );
  NAND2_X2 U2880 ( .A1(decode_regfile_fpregs_6__31_), .A2(n13374), .ZN(n1647)
         );
  NAND2_X2 U2882 ( .A1(decode_regfile_fpregs_6__30_), .A2(n13373), .ZN(n1648)
         );
  NAND2_X2 U2884 ( .A1(decode_regfile_fpregs_6__2_), .A2(n13373), .ZN(n1649)
         );
  NAND2_X2 U2886 ( .A1(decode_regfile_fpregs_6__29_), .A2(n13373), .ZN(n1650)
         );
  NAND2_X2 U2888 ( .A1(decode_regfile_fpregs_6__28_), .A2(n13373), .ZN(n1651)
         );
  NAND2_X2 U2890 ( .A1(decode_regfile_fpregs_6__27_), .A2(n13373), .ZN(n1652)
         );
  NAND2_X2 U2892 ( .A1(decode_regfile_fpregs_6__26_), .A2(n13373), .ZN(n1653)
         );
  NAND2_X2 U2894 ( .A1(decode_regfile_fpregs_6__25_), .A2(n13373), .ZN(n1654)
         );
  NAND2_X2 U2896 ( .A1(decode_regfile_fpregs_6__24_), .A2(n13373), .ZN(n1655)
         );
  NAND2_X2 U2898 ( .A1(decode_regfile_fpregs_6__23_), .A2(n13373), .ZN(n1656)
         );
  NAND2_X2 U2900 ( .A1(decode_regfile_fpregs_6__22_), .A2(n13373), .ZN(n1657)
         );
  NAND2_X2 U2902 ( .A1(decode_regfile_fpregs_6__21_), .A2(n13373), .ZN(n1658)
         );
  NAND2_X2 U2904 ( .A1(decode_regfile_fpregs_6__20_), .A2(n13373), .ZN(n1659)
         );
  NAND2_X2 U2906 ( .A1(decode_regfile_fpregs_6__1_), .A2(n13373), .ZN(n1660)
         );
  NAND2_X2 U2908 ( .A1(decode_regfile_fpregs_6__19_), .A2(n13373), .ZN(n1661)
         );
  NAND2_X2 U2910 ( .A1(decode_regfile_fpregs_6__18_), .A2(n13373), .ZN(n1662)
         );
  NAND2_X2 U2912 ( .A1(decode_regfile_fpregs_6__17_), .A2(n13373), .ZN(n1663)
         );
  NAND2_X2 U2914 ( .A1(decode_regfile_fpregs_6__16_), .A2(n13372), .ZN(n1664)
         );
  NAND2_X2 U2916 ( .A1(decode_regfile_fpregs_6__15_), .A2(n13372), .ZN(n1665)
         );
  NAND2_X2 U2918 ( .A1(decode_regfile_fpregs_6__14_), .A2(n13373), .ZN(n1666)
         );
  NAND2_X2 U2920 ( .A1(decode_regfile_fpregs_6__13_), .A2(n13372), .ZN(n1667)
         );
  NAND2_X2 U2922 ( .A1(decode_regfile_fpregs_6__12_), .A2(n13372), .ZN(n1668)
         );
  NAND2_X2 U2924 ( .A1(decode_regfile_fpregs_6__11_), .A2(n13373), .ZN(n1669)
         );
  NAND2_X2 U2926 ( .A1(decode_regfile_fpregs_6__10_), .A2(n13372), .ZN(n1670)
         );
  NAND2_X2 U2928 ( .A1(decode_regfile_fpregs_6__0_), .A2(n13373), .ZN(n1671)
         );
  NAND2_X2 U2931 ( .A1(decode_regfile_fpregs_5__9_), .A2(n13367), .ZN(n1673)
         );
  NAND2_X2 U2933 ( .A1(decode_regfile_fpregs_5__8_), .A2(n1672), .ZN(n1674) );
  NAND2_X2 U2935 ( .A1(decode_regfile_fpregs_5__7_), .A2(n1672), .ZN(n1675) );
  NAND2_X2 U2937 ( .A1(decode_regfile_fpregs_5__6_), .A2(n1672), .ZN(n1676) );
  NAND2_X2 U2939 ( .A1(decode_regfile_fpregs_5__5_), .A2(n1672), .ZN(n1677) );
  NAND2_X2 U2941 ( .A1(decode_regfile_fpregs_5__4_), .A2(n1672), .ZN(n1678) );
  NAND2_X2 U2943 ( .A1(decode_regfile_fpregs_5__3_), .A2(n1672), .ZN(n1679) );
  NAND2_X2 U2945 ( .A1(decode_regfile_fpregs_5__31_), .A2(n1672), .ZN(n1680)
         );
  NAND2_X2 U2947 ( .A1(decode_regfile_fpregs_5__30_), .A2(n13368), .ZN(n1681)
         );
  NAND2_X2 U2949 ( .A1(decode_regfile_fpregs_5__2_), .A2(n13368), .ZN(n1682)
         );
  NAND2_X2 U2951 ( .A1(decode_regfile_fpregs_5__29_), .A2(n13368), .ZN(n1683)
         );
  NAND2_X2 U2953 ( .A1(decode_regfile_fpregs_5__28_), .A2(n13368), .ZN(n1684)
         );
  NAND2_X2 U2955 ( .A1(decode_regfile_fpregs_5__27_), .A2(n13368), .ZN(n1685)
         );
  NAND2_X2 U2957 ( .A1(decode_regfile_fpregs_5__26_), .A2(n13368), .ZN(n1686)
         );
  NAND2_X2 U2959 ( .A1(decode_regfile_fpregs_5__25_), .A2(n13368), .ZN(n1687)
         );
  NAND2_X2 U2961 ( .A1(decode_regfile_fpregs_5__24_), .A2(n13368), .ZN(n1688)
         );
  NAND2_X2 U2963 ( .A1(decode_regfile_fpregs_5__23_), .A2(n13368), .ZN(n1689)
         );
  NAND2_X2 U2965 ( .A1(decode_regfile_fpregs_5__22_), .A2(n13368), .ZN(n1690)
         );
  NAND2_X2 U2967 ( .A1(decode_regfile_fpregs_5__21_), .A2(n13368), .ZN(n1691)
         );
  NAND2_X2 U2969 ( .A1(decode_regfile_fpregs_5__20_), .A2(n13368), .ZN(n1692)
         );
  NAND2_X2 U2971 ( .A1(decode_regfile_fpregs_5__1_), .A2(n13368), .ZN(n1693)
         );
  NAND2_X2 U2973 ( .A1(decode_regfile_fpregs_5__19_), .A2(n13368), .ZN(n1694)
         );
  NAND2_X2 U2975 ( .A1(decode_regfile_fpregs_5__18_), .A2(n13368), .ZN(n1695)
         );
  NAND2_X2 U2977 ( .A1(decode_regfile_fpregs_5__17_), .A2(n13368), .ZN(n1696)
         );
  NAND2_X2 U2979 ( .A1(decode_regfile_fpregs_5__16_), .A2(n13367), .ZN(n1697)
         );
  NAND2_X2 U2981 ( .A1(decode_regfile_fpregs_5__15_), .A2(n13367), .ZN(n1698)
         );
  NAND2_X2 U2983 ( .A1(decode_regfile_fpregs_5__14_), .A2(n13368), .ZN(n1699)
         );
  NAND2_X2 U2985 ( .A1(decode_regfile_fpregs_5__13_), .A2(n13367), .ZN(n1700)
         );
  NAND2_X2 U2987 ( .A1(decode_regfile_fpregs_5__12_), .A2(n13367), .ZN(n1701)
         );
  NAND2_X2 U2989 ( .A1(decode_regfile_fpregs_5__11_), .A2(n13368), .ZN(n1702)
         );
  NAND2_X2 U2991 ( .A1(decode_regfile_fpregs_5__10_), .A2(n13367), .ZN(n1703)
         );
  NAND2_X2 U2993 ( .A1(decode_regfile_fpregs_5__0_), .A2(n13368), .ZN(n1704)
         );
  NAND2_X2 U2994 ( .A1(n1638), .A2(n800), .ZN(n1672) );
  NAND2_X2 U2996 ( .A1(decode_regfile_fpregs_4__9_), .A2(n13362), .ZN(n1706)
         );
  NAND2_X2 U2998 ( .A1(decode_regfile_fpregs_4__8_), .A2(n1705), .ZN(n1707) );
  NAND2_X2 U3000 ( .A1(decode_regfile_fpregs_4__7_), .A2(n1705), .ZN(n1708) );
  NAND2_X2 U3002 ( .A1(decode_regfile_fpregs_4__6_), .A2(n1705), .ZN(n1709) );
  NAND2_X2 U3004 ( .A1(decode_regfile_fpregs_4__5_), .A2(n1705), .ZN(n1710) );
  NAND2_X2 U3006 ( .A1(decode_regfile_fpregs_4__4_), .A2(n1705), .ZN(n1711) );
  NAND2_X2 U3008 ( .A1(decode_regfile_fpregs_4__3_), .A2(n1705), .ZN(n1712) );
  NAND2_X2 U3010 ( .A1(decode_regfile_fpregs_4__31_), .A2(n1705), .ZN(n1713)
         );
  NAND2_X2 U3012 ( .A1(decode_regfile_fpregs_4__30_), .A2(n13363), .ZN(n1714)
         );
  NAND2_X2 U3014 ( .A1(decode_regfile_fpregs_4__2_), .A2(n13363), .ZN(n1715)
         );
  NAND2_X2 U3016 ( .A1(decode_regfile_fpregs_4__29_), .A2(n13363), .ZN(n1716)
         );
  NAND2_X2 U3018 ( .A1(decode_regfile_fpregs_4__28_), .A2(n13363), .ZN(n1717)
         );
  NAND2_X2 U3020 ( .A1(decode_regfile_fpregs_4__27_), .A2(n13363), .ZN(n1718)
         );
  NAND2_X2 U3022 ( .A1(decode_regfile_fpregs_4__26_), .A2(n13363), .ZN(n1719)
         );
  NAND2_X2 U3024 ( .A1(decode_regfile_fpregs_4__25_), .A2(n13363), .ZN(n1720)
         );
  NAND2_X2 U3026 ( .A1(decode_regfile_fpregs_4__24_), .A2(n13363), .ZN(n1721)
         );
  NAND2_X2 U3028 ( .A1(decode_regfile_fpregs_4__23_), .A2(n13363), .ZN(n1722)
         );
  NAND2_X2 U3030 ( .A1(decode_regfile_fpregs_4__22_), .A2(n13363), .ZN(n1723)
         );
  NAND2_X2 U3032 ( .A1(decode_regfile_fpregs_4__21_), .A2(n13363), .ZN(n1724)
         );
  NAND2_X2 U3034 ( .A1(decode_regfile_fpregs_4__20_), .A2(n13363), .ZN(n1725)
         );
  NAND2_X2 U3036 ( .A1(decode_regfile_fpregs_4__1_), .A2(n13363), .ZN(n1726)
         );
  NAND2_X2 U3038 ( .A1(decode_regfile_fpregs_4__19_), .A2(n13363), .ZN(n1727)
         );
  NAND2_X2 U3040 ( .A1(decode_regfile_fpregs_4__18_), .A2(n13363), .ZN(n1728)
         );
  NAND2_X2 U3042 ( .A1(decode_regfile_fpregs_4__17_), .A2(n13363), .ZN(n1729)
         );
  NAND2_X2 U3044 ( .A1(decode_regfile_fpregs_4__16_), .A2(n13362), .ZN(n1730)
         );
  NAND2_X2 U3046 ( .A1(decode_regfile_fpregs_4__15_), .A2(n13362), .ZN(n1731)
         );
  NAND2_X2 U3048 ( .A1(decode_regfile_fpregs_4__14_), .A2(n13363), .ZN(n1732)
         );
  NAND2_X2 U3050 ( .A1(decode_regfile_fpregs_4__13_), .A2(n13362), .ZN(n1733)
         );
  NAND2_X2 U3052 ( .A1(decode_regfile_fpregs_4__12_), .A2(n13362), .ZN(n1734)
         );
  NAND2_X2 U3054 ( .A1(decode_regfile_fpregs_4__11_), .A2(n13363), .ZN(n1735)
         );
  NAND2_X2 U3056 ( .A1(decode_regfile_fpregs_4__10_), .A2(n13362), .ZN(n1736)
         );
  NAND2_X2 U3058 ( .A1(decode_regfile_fpregs_4__0_), .A2(n13363), .ZN(n1737)
         );
  NAND2_X2 U3059 ( .A1(n1638), .A2(n834), .ZN(n1705) );
  AND2_X2 U3060 ( .A1(n1738), .A2(n530), .ZN(n1638) );
  NAND2_X2 U3062 ( .A1(decode_regfile_fpregs_3__9_), .A2(n13357), .ZN(n1740)
         );
  NAND2_X2 U3064 ( .A1(decode_regfile_fpregs_3__8_), .A2(n13359), .ZN(n1741)
         );
  NAND2_X2 U3066 ( .A1(decode_regfile_fpregs_3__7_), .A2(n13359), .ZN(n1742)
         );
  NAND2_X2 U3068 ( .A1(decode_regfile_fpregs_3__6_), .A2(n13359), .ZN(n1743)
         );
  NAND2_X2 U3070 ( .A1(decode_regfile_fpregs_3__5_), .A2(n13359), .ZN(n1744)
         );
  NAND2_X2 U3072 ( .A1(decode_regfile_fpregs_3__4_), .A2(n13359), .ZN(n1745)
         );
  NAND2_X2 U3074 ( .A1(decode_regfile_fpregs_3__3_), .A2(n13359), .ZN(n1746)
         );
  NAND2_X2 U3076 ( .A1(decode_regfile_fpregs_3__31_), .A2(n13359), .ZN(n1747)
         );
  NAND2_X2 U3078 ( .A1(decode_regfile_fpregs_3__30_), .A2(n13358), .ZN(n1748)
         );
  NAND2_X2 U3080 ( .A1(decode_regfile_fpregs_3__2_), .A2(n13358), .ZN(n1749)
         );
  NAND2_X2 U3082 ( .A1(decode_regfile_fpregs_3__29_), .A2(n13358), .ZN(n1750)
         );
  NAND2_X2 U3084 ( .A1(decode_regfile_fpregs_3__28_), .A2(n13358), .ZN(n1751)
         );
  NAND2_X2 U3086 ( .A1(decode_regfile_fpregs_3__27_), .A2(n13358), .ZN(n1752)
         );
  NAND2_X2 U3088 ( .A1(decode_regfile_fpregs_3__26_), .A2(n13358), .ZN(n1753)
         );
  NAND2_X2 U3090 ( .A1(decode_regfile_fpregs_3__25_), .A2(n13358), .ZN(n1754)
         );
  NAND2_X2 U3092 ( .A1(decode_regfile_fpregs_3__24_), .A2(n13358), .ZN(n1755)
         );
  NAND2_X2 U3094 ( .A1(decode_regfile_fpregs_3__23_), .A2(n13358), .ZN(n1756)
         );
  NAND2_X2 U3096 ( .A1(decode_regfile_fpregs_3__22_), .A2(n13358), .ZN(n1757)
         );
  NAND2_X2 U3098 ( .A1(decode_regfile_fpregs_3__21_), .A2(n13358), .ZN(n1758)
         );
  NAND2_X2 U3100 ( .A1(decode_regfile_fpregs_3__20_), .A2(n13358), .ZN(n1759)
         );
  NAND2_X2 U3102 ( .A1(decode_regfile_fpregs_3__1_), .A2(n13358), .ZN(n1760)
         );
  NAND2_X2 U3104 ( .A1(decode_regfile_fpregs_3__19_), .A2(n13358), .ZN(n1761)
         );
  NAND2_X2 U3106 ( .A1(decode_regfile_fpregs_3__18_), .A2(n13358), .ZN(n1762)
         );
  NAND2_X2 U3108 ( .A1(decode_regfile_fpregs_3__17_), .A2(n13358), .ZN(n1763)
         );
  NAND2_X2 U3110 ( .A1(decode_regfile_fpregs_3__16_), .A2(n13357), .ZN(n1764)
         );
  NAND2_X2 U3112 ( .A1(decode_regfile_fpregs_3__15_), .A2(n13357), .ZN(n1765)
         );
  NAND2_X2 U3114 ( .A1(decode_regfile_fpregs_3__14_), .A2(n13358), .ZN(n1766)
         );
  NAND2_X2 U3116 ( .A1(decode_regfile_fpregs_3__13_), .A2(n13357), .ZN(n1767)
         );
  NAND2_X2 U3118 ( .A1(decode_regfile_fpregs_3__12_), .A2(n13357), .ZN(n1768)
         );
  NAND2_X2 U3120 ( .A1(decode_regfile_fpregs_3__11_), .A2(n13358), .ZN(n1769)
         );
  NAND2_X2 U3122 ( .A1(decode_regfile_fpregs_3__10_), .A2(n13357), .ZN(n1770)
         );
  NAND2_X2 U3124 ( .A1(decode_regfile_fpregs_3__0_), .A2(n13358), .ZN(n1771)
         );
  NAND2_X2 U3127 ( .A1(decode_regfile_fpregs_31__9_), .A2(n13352), .ZN(n1774)
         );
  NAND2_X2 U3129 ( .A1(decode_regfile_fpregs_31__8_), .A2(n13354), .ZN(n1775)
         );
  NAND2_X2 U3131 ( .A1(decode_regfile_fpregs_31__7_), .A2(n13354), .ZN(n1776)
         );
  NAND2_X2 U3133 ( .A1(decode_regfile_fpregs_31__6_), .A2(n13354), .ZN(n1777)
         );
  NAND2_X2 U3135 ( .A1(decode_regfile_fpregs_31__5_), .A2(n13354), .ZN(n1778)
         );
  NAND2_X2 U3137 ( .A1(decode_regfile_fpregs_31__4_), .A2(n13354), .ZN(n1779)
         );
  NAND2_X2 U3139 ( .A1(decode_regfile_fpregs_31__3_), .A2(n13354), .ZN(n1780)
         );
  NAND2_X2 U3141 ( .A1(decode_regfile_fpregs_31__31_), .A2(n13354), .ZN(n1781)
         );
  NAND2_X2 U3143 ( .A1(decode_regfile_fpregs_31__30_), .A2(n13353), .ZN(n1782)
         );
  NAND2_X2 U3145 ( .A1(decode_regfile_fpregs_31__2_), .A2(n13353), .ZN(n1783)
         );
  NAND2_X2 U3147 ( .A1(decode_regfile_fpregs_31__29_), .A2(n13353), .ZN(n1784)
         );
  NAND2_X2 U3149 ( .A1(decode_regfile_fpregs_31__28_), .A2(n13353), .ZN(n1785)
         );
  NAND2_X2 U3151 ( .A1(decode_regfile_fpregs_31__27_), .A2(n13353), .ZN(n1786)
         );
  NAND2_X2 U3153 ( .A1(decode_regfile_fpregs_31__26_), .A2(n13353), .ZN(n1787)
         );
  NAND2_X2 U3155 ( .A1(decode_regfile_fpregs_31__25_), .A2(n13353), .ZN(n1788)
         );
  NAND2_X2 U3157 ( .A1(decode_regfile_fpregs_31__24_), .A2(n13353), .ZN(n1789)
         );
  NAND2_X2 U3159 ( .A1(decode_regfile_fpregs_31__23_), .A2(n13353), .ZN(n1790)
         );
  NAND2_X2 U3161 ( .A1(decode_regfile_fpregs_31__22_), .A2(n13353), .ZN(n1791)
         );
  NAND2_X2 U3163 ( .A1(decode_regfile_fpregs_31__21_), .A2(n13353), .ZN(n1792)
         );
  NAND2_X2 U3165 ( .A1(decode_regfile_fpregs_31__20_), .A2(n13353), .ZN(n1793)
         );
  NAND2_X2 U3167 ( .A1(decode_regfile_fpregs_31__1_), .A2(n13353), .ZN(n1794)
         );
  NAND2_X2 U3169 ( .A1(decode_regfile_fpregs_31__19_), .A2(n13353), .ZN(n1795)
         );
  NAND2_X2 U3171 ( .A1(decode_regfile_fpregs_31__18_), .A2(n13353), .ZN(n1796)
         );
  NAND2_X2 U3173 ( .A1(decode_regfile_fpregs_31__17_), .A2(n13353), .ZN(n1797)
         );
  NAND2_X2 U3175 ( .A1(decode_regfile_fpregs_31__16_), .A2(n13352), .ZN(n1798)
         );
  NAND2_X2 U3177 ( .A1(decode_regfile_fpregs_31__15_), .A2(n13352), .ZN(n1799)
         );
  NAND2_X2 U3179 ( .A1(decode_regfile_fpregs_31__14_), .A2(n13353), .ZN(n1800)
         );
  NAND2_X2 U3181 ( .A1(decode_regfile_fpregs_31__13_), .A2(n13352), .ZN(n1801)
         );
  NAND2_X2 U3183 ( .A1(decode_regfile_fpregs_31__12_), .A2(n13352), .ZN(n1802)
         );
  NAND2_X2 U3185 ( .A1(decode_regfile_fpregs_31__11_), .A2(n13353), .ZN(n1803)
         );
  NAND2_X2 U3187 ( .A1(decode_regfile_fpregs_31__10_), .A2(n13352), .ZN(n1804)
         );
  NAND2_X2 U3189 ( .A1(decode_regfile_fpregs_31__0_), .A2(n13353), .ZN(n1805)
         );
  NAND2_X2 U3192 ( .A1(decode_regfile_fpregs_30__9_), .A2(n13347), .ZN(n1808)
         );
  NAND2_X2 U3194 ( .A1(decode_regfile_fpregs_30__8_), .A2(n13349), .ZN(n1809)
         );
  NAND2_X2 U3196 ( .A1(decode_regfile_fpregs_30__7_), .A2(n13349), .ZN(n1810)
         );
  NAND2_X2 U3198 ( .A1(decode_regfile_fpregs_30__6_), .A2(n13349), .ZN(n1811)
         );
  NAND2_X2 U3200 ( .A1(decode_regfile_fpregs_30__5_), .A2(n13349), .ZN(n1812)
         );
  NAND2_X2 U3202 ( .A1(decode_regfile_fpregs_30__4_), .A2(n13349), .ZN(n1813)
         );
  NAND2_X2 U3204 ( .A1(decode_regfile_fpregs_30__3_), .A2(n13349), .ZN(n1814)
         );
  NAND2_X2 U3206 ( .A1(decode_regfile_fpregs_30__31_), .A2(n13349), .ZN(n1815)
         );
  NAND2_X2 U3208 ( .A1(decode_regfile_fpregs_30__30_), .A2(n13348), .ZN(n1816)
         );
  NAND2_X2 U3210 ( .A1(decode_regfile_fpregs_30__2_), .A2(n13348), .ZN(n1817)
         );
  NAND2_X2 U3212 ( .A1(decode_regfile_fpregs_30__29_), .A2(n13348), .ZN(n1818)
         );
  NAND2_X2 U3214 ( .A1(decode_regfile_fpregs_30__28_), .A2(n13348), .ZN(n1819)
         );
  NAND2_X2 U3216 ( .A1(decode_regfile_fpregs_30__27_), .A2(n13348), .ZN(n1820)
         );
  NAND2_X2 U3218 ( .A1(decode_regfile_fpregs_30__26_), .A2(n13348), .ZN(n1821)
         );
  NAND2_X2 U3220 ( .A1(decode_regfile_fpregs_30__25_), .A2(n13348), .ZN(n1822)
         );
  NAND2_X2 U3222 ( .A1(decode_regfile_fpregs_30__24_), .A2(n13348), .ZN(n1823)
         );
  NAND2_X2 U3224 ( .A1(decode_regfile_fpregs_30__23_), .A2(n13348), .ZN(n1824)
         );
  NAND2_X2 U3226 ( .A1(decode_regfile_fpregs_30__22_), .A2(n13348), .ZN(n1825)
         );
  NAND2_X2 U3228 ( .A1(decode_regfile_fpregs_30__21_), .A2(n13348), .ZN(n1826)
         );
  NAND2_X2 U3230 ( .A1(decode_regfile_fpregs_30__20_), .A2(n13348), .ZN(n1827)
         );
  NAND2_X2 U3232 ( .A1(decode_regfile_fpregs_30__1_), .A2(n13348), .ZN(n1828)
         );
  NAND2_X2 U3234 ( .A1(decode_regfile_fpregs_30__19_), .A2(n13348), .ZN(n1829)
         );
  NAND2_X2 U3236 ( .A1(decode_regfile_fpregs_30__18_), .A2(n13348), .ZN(n1830)
         );
  NAND2_X2 U3238 ( .A1(decode_regfile_fpregs_30__17_), .A2(n13348), .ZN(n1831)
         );
  NAND2_X2 U3240 ( .A1(decode_regfile_fpregs_30__16_), .A2(n13347), .ZN(n1832)
         );
  NAND2_X2 U3242 ( .A1(decode_regfile_fpregs_30__15_), .A2(n13347), .ZN(n1833)
         );
  NAND2_X2 U3244 ( .A1(decode_regfile_fpregs_30__14_), .A2(n13348), .ZN(n1834)
         );
  NAND2_X2 U3246 ( .A1(decode_regfile_fpregs_30__13_), .A2(n13347), .ZN(n1835)
         );
  NAND2_X2 U3248 ( .A1(decode_regfile_fpregs_30__12_), .A2(n13347), .ZN(n1836)
         );
  NAND2_X2 U3250 ( .A1(decode_regfile_fpregs_30__11_), .A2(n13348), .ZN(n1837)
         );
  NAND2_X2 U3252 ( .A1(decode_regfile_fpregs_30__10_), .A2(n13347), .ZN(n1838)
         );
  NAND2_X2 U3254 ( .A1(decode_regfile_fpregs_30__0_), .A2(n13348), .ZN(n1839)
         );
  NAND2_X2 U3257 ( .A1(decode_regfile_fpregs_2__9_), .A2(n13342), .ZN(n1841)
         );
  NAND2_X2 U3259 ( .A1(decode_regfile_fpregs_2__8_), .A2(n13344), .ZN(n1842)
         );
  NAND2_X2 U3261 ( .A1(decode_regfile_fpregs_2__7_), .A2(n13344), .ZN(n1843)
         );
  NAND2_X2 U3263 ( .A1(decode_regfile_fpregs_2__6_), .A2(n13344), .ZN(n1844)
         );
  NAND2_X2 U3265 ( .A1(decode_regfile_fpregs_2__5_), .A2(n13344), .ZN(n1845)
         );
  NAND2_X2 U3267 ( .A1(decode_regfile_fpregs_2__4_), .A2(n13344), .ZN(n1846)
         );
  NAND2_X2 U3269 ( .A1(decode_regfile_fpregs_2__3_), .A2(n13344), .ZN(n1847)
         );
  NAND2_X2 U3271 ( .A1(decode_regfile_fpregs_2__31_), .A2(n13344), .ZN(n1848)
         );
  NAND2_X2 U3273 ( .A1(decode_regfile_fpregs_2__30_), .A2(n13343), .ZN(n1849)
         );
  NAND2_X2 U3275 ( .A1(decode_regfile_fpregs_2__2_), .A2(n13343), .ZN(n1850)
         );
  NAND2_X2 U3277 ( .A1(decode_regfile_fpregs_2__29_), .A2(n13343), .ZN(n1851)
         );
  NAND2_X2 U3279 ( .A1(decode_regfile_fpregs_2__28_), .A2(n13343), .ZN(n1852)
         );
  NAND2_X2 U3281 ( .A1(decode_regfile_fpregs_2__27_), .A2(n13343), .ZN(n1853)
         );
  NAND2_X2 U3283 ( .A1(decode_regfile_fpregs_2__26_), .A2(n13343), .ZN(n1854)
         );
  NAND2_X2 U3285 ( .A1(decode_regfile_fpregs_2__25_), .A2(n13343), .ZN(n1855)
         );
  NAND2_X2 U3287 ( .A1(decode_regfile_fpregs_2__24_), .A2(n13343), .ZN(n1856)
         );
  NAND2_X2 U3289 ( .A1(decode_regfile_fpregs_2__23_), .A2(n13343), .ZN(n1857)
         );
  NAND2_X2 U3291 ( .A1(decode_regfile_fpregs_2__22_), .A2(n13343), .ZN(n1858)
         );
  NAND2_X2 U3293 ( .A1(decode_regfile_fpregs_2__21_), .A2(n13343), .ZN(n1859)
         );
  NAND2_X2 U3295 ( .A1(decode_regfile_fpregs_2__20_), .A2(n13343), .ZN(n1860)
         );
  NAND2_X2 U3297 ( .A1(decode_regfile_fpregs_2__1_), .A2(n13343), .ZN(n1861)
         );
  NAND2_X2 U3299 ( .A1(decode_regfile_fpregs_2__19_), .A2(n13343), .ZN(n1862)
         );
  NAND2_X2 U3301 ( .A1(decode_regfile_fpregs_2__18_), .A2(n13343), .ZN(n1863)
         );
  NAND2_X2 U3303 ( .A1(decode_regfile_fpregs_2__17_), .A2(n13343), .ZN(n1864)
         );
  NAND2_X2 U3305 ( .A1(decode_regfile_fpregs_2__16_), .A2(n13342), .ZN(n1865)
         );
  NAND2_X2 U3307 ( .A1(decode_regfile_fpregs_2__15_), .A2(n13342), .ZN(n1866)
         );
  NAND2_X2 U3309 ( .A1(decode_regfile_fpregs_2__14_), .A2(n13343), .ZN(n1867)
         );
  NAND2_X2 U3311 ( .A1(decode_regfile_fpregs_2__13_), .A2(n13342), .ZN(n1868)
         );
  NAND2_X2 U3313 ( .A1(decode_regfile_fpregs_2__12_), .A2(n13342), .ZN(n1869)
         );
  NAND2_X2 U3315 ( .A1(decode_regfile_fpregs_2__11_), .A2(n13343), .ZN(n1870)
         );
  NAND2_X2 U3317 ( .A1(decode_regfile_fpregs_2__10_), .A2(n13342), .ZN(n1871)
         );
  NAND2_X2 U3319 ( .A1(decode_regfile_fpregs_2__0_), .A2(n13343), .ZN(n1872)
         );
  NAND2_X2 U3322 ( .A1(decode_regfile_fpregs_29__9_), .A2(n13337), .ZN(n1874)
         );
  NAND2_X2 U3324 ( .A1(decode_regfile_fpregs_29__8_), .A2(n1873), .ZN(n1875)
         );
  NAND2_X2 U3326 ( .A1(decode_regfile_fpregs_29__7_), .A2(n1873), .ZN(n1876)
         );
  NAND2_X2 U3328 ( .A1(decode_regfile_fpregs_29__6_), .A2(n1873), .ZN(n1877)
         );
  NAND2_X2 U3330 ( .A1(decode_regfile_fpregs_29__5_), .A2(n1873), .ZN(n1878)
         );
  NAND2_X2 U3332 ( .A1(decode_regfile_fpregs_29__4_), .A2(n1873), .ZN(n1879)
         );
  NAND2_X2 U3334 ( .A1(decode_regfile_fpregs_29__3_), .A2(n1873), .ZN(n1880)
         );
  NAND2_X2 U3336 ( .A1(decode_regfile_fpregs_29__31_), .A2(n1873), .ZN(n1881)
         );
  NAND2_X2 U3338 ( .A1(decode_regfile_fpregs_29__30_), .A2(n13338), .ZN(n1882)
         );
  NAND2_X2 U3340 ( .A1(decode_regfile_fpregs_29__2_), .A2(n13338), .ZN(n1883)
         );
  NAND2_X2 U3342 ( .A1(decode_regfile_fpregs_29__29_), .A2(n13338), .ZN(n1884)
         );
  NAND2_X2 U3344 ( .A1(decode_regfile_fpregs_29__28_), .A2(n13338), .ZN(n1885)
         );
  NAND2_X2 U3346 ( .A1(decode_regfile_fpregs_29__27_), .A2(n13338), .ZN(n1886)
         );
  NAND2_X2 U3348 ( .A1(decode_regfile_fpregs_29__26_), .A2(n13338), .ZN(n1887)
         );
  NAND2_X2 U3350 ( .A1(decode_regfile_fpregs_29__25_), .A2(n13338), .ZN(n1888)
         );
  NAND2_X2 U3352 ( .A1(decode_regfile_fpregs_29__24_), .A2(n13338), .ZN(n1889)
         );
  NAND2_X2 U3354 ( .A1(decode_regfile_fpregs_29__23_), .A2(n13338), .ZN(n1890)
         );
  NAND2_X2 U3356 ( .A1(decode_regfile_fpregs_29__22_), .A2(n13338), .ZN(n1891)
         );
  NAND2_X2 U3358 ( .A1(decode_regfile_fpregs_29__21_), .A2(n13338), .ZN(n1892)
         );
  NAND2_X2 U3360 ( .A1(decode_regfile_fpregs_29__20_), .A2(n13338), .ZN(n1893)
         );
  NAND2_X2 U3362 ( .A1(decode_regfile_fpregs_29__1_), .A2(n13338), .ZN(n1894)
         );
  NAND2_X2 U3364 ( .A1(decode_regfile_fpregs_29__19_), .A2(n13338), .ZN(n1895)
         );
  NAND2_X2 U3366 ( .A1(decode_regfile_fpregs_29__18_), .A2(n13338), .ZN(n1896)
         );
  NAND2_X2 U3368 ( .A1(decode_regfile_fpregs_29__17_), .A2(n13338), .ZN(n1897)
         );
  NAND2_X2 U3370 ( .A1(decode_regfile_fpregs_29__16_), .A2(n13337), .ZN(n1898)
         );
  NAND2_X2 U3372 ( .A1(decode_regfile_fpregs_29__15_), .A2(n13337), .ZN(n1899)
         );
  NAND2_X2 U3374 ( .A1(decode_regfile_fpregs_29__14_), .A2(n13338), .ZN(n1900)
         );
  NAND2_X2 U3376 ( .A1(decode_regfile_fpregs_29__13_), .A2(n13337), .ZN(n1901)
         );
  NAND2_X2 U3378 ( .A1(decode_regfile_fpregs_29__12_), .A2(n13337), .ZN(n1902)
         );
  NAND2_X2 U3380 ( .A1(decode_regfile_fpregs_29__11_), .A2(n13338), .ZN(n1903)
         );
  NAND2_X2 U3382 ( .A1(decode_regfile_fpregs_29__10_), .A2(n13337), .ZN(n1904)
         );
  NAND2_X2 U3384 ( .A1(decode_regfile_fpregs_29__0_), .A2(n13338), .ZN(n1905)
         );
  NAND2_X2 U3385 ( .A1(n1806), .A2(n800), .ZN(n1873) );
  NAND2_X2 U3387 ( .A1(decode_regfile_fpregs_28__9_), .A2(n13332), .ZN(n1907)
         );
  NAND2_X2 U3389 ( .A1(decode_regfile_fpregs_28__8_), .A2(n1906), .ZN(n1908)
         );
  NAND2_X2 U3391 ( .A1(decode_regfile_fpregs_28__7_), .A2(n1906), .ZN(n1909)
         );
  NAND2_X2 U3393 ( .A1(decode_regfile_fpregs_28__6_), .A2(n1906), .ZN(n1910)
         );
  NAND2_X2 U3395 ( .A1(decode_regfile_fpregs_28__5_), .A2(n1906), .ZN(n1911)
         );
  NAND2_X2 U3397 ( .A1(decode_regfile_fpregs_28__4_), .A2(n1906), .ZN(n1912)
         );
  NAND2_X2 U3399 ( .A1(decode_regfile_fpregs_28__3_), .A2(n1906), .ZN(n1913)
         );
  NAND2_X2 U3401 ( .A1(decode_regfile_fpregs_28__31_), .A2(n1906), .ZN(n1914)
         );
  NAND2_X2 U3403 ( .A1(decode_regfile_fpregs_28__30_), .A2(n13333), .ZN(n1915)
         );
  NAND2_X2 U3405 ( .A1(decode_regfile_fpregs_28__2_), .A2(n13333), .ZN(n1916)
         );
  NAND2_X2 U3407 ( .A1(decode_regfile_fpregs_28__29_), .A2(n13333), .ZN(n1917)
         );
  NAND2_X2 U3409 ( .A1(decode_regfile_fpregs_28__28_), .A2(n13333), .ZN(n1918)
         );
  NAND2_X2 U3411 ( .A1(decode_regfile_fpregs_28__27_), .A2(n13333), .ZN(n1919)
         );
  NAND2_X2 U3413 ( .A1(decode_regfile_fpregs_28__26_), .A2(n13333), .ZN(n1920)
         );
  NAND2_X2 U3415 ( .A1(decode_regfile_fpregs_28__25_), .A2(n13333), .ZN(n1921)
         );
  NAND2_X2 U3417 ( .A1(decode_regfile_fpregs_28__24_), .A2(n13333), .ZN(n1922)
         );
  NAND2_X2 U3419 ( .A1(decode_regfile_fpregs_28__23_), .A2(n13333), .ZN(n1923)
         );
  NAND2_X2 U3421 ( .A1(decode_regfile_fpregs_28__22_), .A2(n13333), .ZN(n1924)
         );
  NAND2_X2 U3423 ( .A1(decode_regfile_fpregs_28__21_), .A2(n13333), .ZN(n1925)
         );
  NAND2_X2 U3425 ( .A1(decode_regfile_fpregs_28__20_), .A2(n13333), .ZN(n1926)
         );
  NAND2_X2 U3427 ( .A1(decode_regfile_fpregs_28__1_), .A2(n13333), .ZN(n1927)
         );
  NAND2_X2 U3429 ( .A1(decode_regfile_fpregs_28__19_), .A2(n13333), .ZN(n1928)
         );
  NAND2_X2 U3431 ( .A1(decode_regfile_fpregs_28__18_), .A2(n13333), .ZN(n1929)
         );
  NAND2_X2 U3433 ( .A1(decode_regfile_fpregs_28__17_), .A2(n13333), .ZN(n1930)
         );
  NAND2_X2 U3435 ( .A1(decode_regfile_fpregs_28__16_), .A2(n13332), .ZN(n1931)
         );
  NAND2_X2 U3437 ( .A1(decode_regfile_fpregs_28__15_), .A2(n13332), .ZN(n1932)
         );
  NAND2_X2 U3439 ( .A1(decode_regfile_fpregs_28__14_), .A2(n13333), .ZN(n1933)
         );
  NAND2_X2 U3441 ( .A1(decode_regfile_fpregs_28__13_), .A2(n13332), .ZN(n1934)
         );
  NAND2_X2 U3443 ( .A1(decode_regfile_fpregs_28__12_), .A2(n13332), .ZN(n1935)
         );
  NAND2_X2 U3445 ( .A1(decode_regfile_fpregs_28__11_), .A2(n13333), .ZN(n1936)
         );
  NAND2_X2 U3447 ( .A1(decode_regfile_fpregs_28__10_), .A2(n13332), .ZN(n1937)
         );
  NAND2_X2 U3449 ( .A1(decode_regfile_fpregs_28__0_), .A2(n13333), .ZN(n1938)
         );
  NAND2_X2 U3450 ( .A1(n1806), .A2(n834), .ZN(n1906) );
  AND2_X2 U3451 ( .A1(n1939), .A2(n836), .ZN(n1806) );
  NAND2_X2 U3453 ( .A1(decode_regfile_fpregs_27__9_), .A2(n13327), .ZN(n1941)
         );
  NAND2_X2 U3455 ( .A1(decode_regfile_fpregs_27__8_), .A2(n13329), .ZN(n1942)
         );
  NAND2_X2 U3457 ( .A1(decode_regfile_fpregs_27__7_), .A2(n13329), .ZN(n1943)
         );
  NAND2_X2 U3459 ( .A1(decode_regfile_fpregs_27__6_), .A2(n13329), .ZN(n1944)
         );
  NAND2_X2 U3461 ( .A1(decode_regfile_fpregs_27__5_), .A2(n13329), .ZN(n1945)
         );
  NAND2_X2 U3463 ( .A1(decode_regfile_fpregs_27__4_), .A2(n13329), .ZN(n1946)
         );
  NAND2_X2 U3465 ( .A1(decode_regfile_fpregs_27__3_), .A2(n13329), .ZN(n1947)
         );
  NAND2_X2 U3467 ( .A1(decode_regfile_fpregs_27__31_), .A2(n13329), .ZN(n1948)
         );
  NAND2_X2 U3469 ( .A1(decode_regfile_fpregs_27__30_), .A2(n13328), .ZN(n1949)
         );
  NAND2_X2 U3471 ( .A1(decode_regfile_fpregs_27__2_), .A2(n13328), .ZN(n1950)
         );
  NAND2_X2 U3473 ( .A1(decode_regfile_fpregs_27__29_), .A2(n13328), .ZN(n1951)
         );
  NAND2_X2 U3475 ( .A1(decode_regfile_fpregs_27__28_), .A2(n13328), .ZN(n1952)
         );
  NAND2_X2 U3477 ( .A1(decode_regfile_fpregs_27__27_), .A2(n13328), .ZN(n1953)
         );
  NAND2_X2 U3479 ( .A1(decode_regfile_fpregs_27__26_), .A2(n13328), .ZN(n1954)
         );
  NAND2_X2 U3481 ( .A1(decode_regfile_fpregs_27__25_), .A2(n13328), .ZN(n1955)
         );
  NAND2_X2 U3483 ( .A1(decode_regfile_fpregs_27__24_), .A2(n13328), .ZN(n1956)
         );
  NAND2_X2 U3485 ( .A1(decode_regfile_fpregs_27__23_), .A2(n13328), .ZN(n1957)
         );
  NAND2_X2 U3487 ( .A1(decode_regfile_fpregs_27__22_), .A2(n13328), .ZN(n1958)
         );
  NAND2_X2 U3489 ( .A1(decode_regfile_fpregs_27__21_), .A2(n13328), .ZN(n1959)
         );
  NAND2_X2 U3491 ( .A1(decode_regfile_fpregs_27__20_), .A2(n13328), .ZN(n1960)
         );
  NAND2_X2 U3493 ( .A1(decode_regfile_fpregs_27__1_), .A2(n13328), .ZN(n1961)
         );
  NAND2_X2 U3495 ( .A1(decode_regfile_fpregs_27__19_), .A2(n13328), .ZN(n1962)
         );
  NAND2_X2 U3497 ( .A1(decode_regfile_fpregs_27__18_), .A2(n13328), .ZN(n1963)
         );
  NAND2_X2 U3499 ( .A1(decode_regfile_fpregs_27__17_), .A2(n13328), .ZN(n1964)
         );
  NAND2_X2 U3501 ( .A1(decode_regfile_fpregs_27__16_), .A2(n13327), .ZN(n1965)
         );
  NAND2_X2 U3503 ( .A1(decode_regfile_fpregs_27__15_), .A2(n13327), .ZN(n1966)
         );
  NAND2_X2 U3505 ( .A1(decode_regfile_fpregs_27__14_), .A2(n13328), .ZN(n1967)
         );
  NAND2_X2 U3507 ( .A1(decode_regfile_fpregs_27__13_), .A2(n13327), .ZN(n1968)
         );
  NAND2_X2 U3509 ( .A1(decode_regfile_fpregs_27__12_), .A2(n13327), .ZN(n1969)
         );
  NAND2_X2 U3511 ( .A1(decode_regfile_fpregs_27__11_), .A2(n13328), .ZN(n1970)
         );
  NAND2_X2 U3513 ( .A1(decode_regfile_fpregs_27__10_), .A2(n13327), .ZN(n1971)
         );
  NAND2_X2 U3515 ( .A1(decode_regfile_fpregs_27__0_), .A2(n13328), .ZN(n1972)
         );
  NAND2_X2 U3518 ( .A1(decode_regfile_fpregs_26__9_), .A2(n13322), .ZN(n1975)
         );
  NAND2_X2 U3520 ( .A1(decode_regfile_fpregs_26__8_), .A2(n13324), .ZN(n1976)
         );
  NAND2_X2 U3522 ( .A1(decode_regfile_fpregs_26__7_), .A2(n13324), .ZN(n1977)
         );
  NAND2_X2 U3524 ( .A1(decode_regfile_fpregs_26__6_), .A2(n13324), .ZN(n1978)
         );
  NAND2_X2 U3526 ( .A1(decode_regfile_fpregs_26__5_), .A2(n13324), .ZN(n1979)
         );
  NAND2_X2 U3528 ( .A1(decode_regfile_fpregs_26__4_), .A2(n13324), .ZN(n1980)
         );
  NAND2_X2 U3530 ( .A1(decode_regfile_fpregs_26__3_), .A2(n13324), .ZN(n1981)
         );
  NAND2_X2 U3532 ( .A1(decode_regfile_fpregs_26__31_), .A2(n13324), .ZN(n1982)
         );
  NAND2_X2 U3534 ( .A1(decode_regfile_fpregs_26__30_), .A2(n13323), .ZN(n1983)
         );
  NAND2_X2 U3536 ( .A1(decode_regfile_fpregs_26__2_), .A2(n13323), .ZN(n1984)
         );
  NAND2_X2 U3538 ( .A1(decode_regfile_fpregs_26__29_), .A2(n13323), .ZN(n1985)
         );
  NAND2_X2 U3540 ( .A1(decode_regfile_fpregs_26__28_), .A2(n13323), .ZN(n1986)
         );
  NAND2_X2 U3542 ( .A1(decode_regfile_fpregs_26__27_), .A2(n13323), .ZN(n1987)
         );
  NAND2_X2 U3544 ( .A1(decode_regfile_fpregs_26__26_), .A2(n13323), .ZN(n1988)
         );
  NAND2_X2 U3546 ( .A1(decode_regfile_fpregs_26__25_), .A2(n13323), .ZN(n1989)
         );
  NAND2_X2 U3548 ( .A1(decode_regfile_fpregs_26__24_), .A2(n13323), .ZN(n1990)
         );
  NAND2_X2 U3550 ( .A1(decode_regfile_fpregs_26__23_), .A2(n13323), .ZN(n1991)
         );
  NAND2_X2 U3552 ( .A1(decode_regfile_fpregs_26__22_), .A2(n13323), .ZN(n1992)
         );
  NAND2_X2 U3554 ( .A1(decode_regfile_fpregs_26__21_), .A2(n13323), .ZN(n1993)
         );
  NAND2_X2 U3556 ( .A1(decode_regfile_fpregs_26__20_), .A2(n13323), .ZN(n1994)
         );
  NAND2_X2 U3558 ( .A1(decode_regfile_fpregs_26__1_), .A2(n13323), .ZN(n1995)
         );
  NAND2_X2 U3560 ( .A1(decode_regfile_fpregs_26__19_), .A2(n13323), .ZN(n1996)
         );
  NAND2_X2 U3562 ( .A1(decode_regfile_fpregs_26__18_), .A2(n13323), .ZN(n1997)
         );
  NAND2_X2 U3564 ( .A1(decode_regfile_fpregs_26__17_), .A2(n13323), .ZN(n1998)
         );
  NAND2_X2 U3566 ( .A1(decode_regfile_fpregs_26__16_), .A2(n13322), .ZN(n1999)
         );
  NAND2_X2 U3568 ( .A1(decode_regfile_fpregs_26__15_), .A2(n13322), .ZN(n2000)
         );
  NAND2_X2 U3570 ( .A1(decode_regfile_fpregs_26__14_), .A2(n13323), .ZN(n2001)
         );
  NAND2_X2 U3572 ( .A1(decode_regfile_fpregs_26__13_), .A2(n13322), .ZN(n2002)
         );
  NAND2_X2 U3574 ( .A1(decode_regfile_fpregs_26__12_), .A2(n13322), .ZN(n2003)
         );
  NAND2_X2 U3576 ( .A1(decode_regfile_fpregs_26__11_), .A2(n13323), .ZN(n2004)
         );
  NAND2_X2 U3578 ( .A1(decode_regfile_fpregs_26__10_), .A2(n13322), .ZN(n2005)
         );
  NAND2_X2 U3580 ( .A1(decode_regfile_fpregs_26__0_), .A2(n13323), .ZN(n2006)
         );
  NAND2_X2 U3583 ( .A1(decode_regfile_fpregs_25__9_), .A2(n13317), .ZN(n2008)
         );
  NAND2_X2 U3585 ( .A1(decode_regfile_fpregs_25__8_), .A2(n2007), .ZN(n2009)
         );
  NAND2_X2 U3587 ( .A1(decode_regfile_fpregs_25__7_), .A2(n2007), .ZN(n2010)
         );
  NAND2_X2 U3589 ( .A1(decode_regfile_fpregs_25__6_), .A2(n2007), .ZN(n2011)
         );
  NAND2_X2 U3591 ( .A1(decode_regfile_fpregs_25__5_), .A2(n2007), .ZN(n2012)
         );
  NAND2_X2 U3593 ( .A1(decode_regfile_fpregs_25__4_), .A2(n2007), .ZN(n2013)
         );
  NAND2_X2 U3595 ( .A1(decode_regfile_fpregs_25__3_), .A2(n2007), .ZN(n2014)
         );
  NAND2_X2 U3597 ( .A1(decode_regfile_fpregs_25__31_), .A2(n2007), .ZN(n2015)
         );
  NAND2_X2 U3599 ( .A1(decode_regfile_fpregs_25__30_), .A2(n13318), .ZN(n2016)
         );
  NAND2_X2 U3601 ( .A1(decode_regfile_fpregs_25__2_), .A2(n13318), .ZN(n2017)
         );
  NAND2_X2 U3603 ( .A1(decode_regfile_fpregs_25__29_), .A2(n13318), .ZN(n2018)
         );
  NAND2_X2 U3605 ( .A1(decode_regfile_fpregs_25__28_), .A2(n13318), .ZN(n2019)
         );
  NAND2_X2 U3607 ( .A1(decode_regfile_fpregs_25__27_), .A2(n13318), .ZN(n2020)
         );
  NAND2_X2 U3609 ( .A1(decode_regfile_fpregs_25__26_), .A2(n13318), .ZN(n2021)
         );
  NAND2_X2 U3611 ( .A1(decode_regfile_fpregs_25__25_), .A2(n13318), .ZN(n2022)
         );
  NAND2_X2 U3613 ( .A1(decode_regfile_fpregs_25__24_), .A2(n13318), .ZN(n2023)
         );
  NAND2_X2 U3615 ( .A1(decode_regfile_fpregs_25__23_), .A2(n13318), .ZN(n2024)
         );
  NAND2_X2 U3617 ( .A1(decode_regfile_fpregs_25__22_), .A2(n13318), .ZN(n2025)
         );
  NAND2_X2 U3619 ( .A1(decode_regfile_fpregs_25__21_), .A2(n13318), .ZN(n2026)
         );
  NAND2_X2 U3621 ( .A1(decode_regfile_fpregs_25__20_), .A2(n13318), .ZN(n2027)
         );
  NAND2_X2 U3623 ( .A1(decode_regfile_fpregs_25__1_), .A2(n13318), .ZN(n2028)
         );
  NAND2_X2 U3625 ( .A1(decode_regfile_fpregs_25__19_), .A2(n13318), .ZN(n2029)
         );
  NAND2_X2 U3627 ( .A1(decode_regfile_fpregs_25__18_), .A2(n13318), .ZN(n2030)
         );
  NAND2_X2 U3629 ( .A1(decode_regfile_fpregs_25__17_), .A2(n13318), .ZN(n2031)
         );
  NAND2_X2 U3631 ( .A1(decode_regfile_fpregs_25__16_), .A2(n13317), .ZN(n2032)
         );
  NAND2_X2 U3633 ( .A1(decode_regfile_fpregs_25__15_), .A2(n13317), .ZN(n2033)
         );
  NAND2_X2 U3635 ( .A1(decode_regfile_fpregs_25__14_), .A2(n13318), .ZN(n2034)
         );
  NAND2_X2 U3637 ( .A1(decode_regfile_fpregs_25__13_), .A2(n13317), .ZN(n2035)
         );
  NAND2_X2 U3639 ( .A1(decode_regfile_fpregs_25__12_), .A2(n13317), .ZN(n2036)
         );
  NAND2_X2 U3641 ( .A1(decode_regfile_fpregs_25__11_), .A2(n13318), .ZN(n2037)
         );
  NAND2_X2 U3643 ( .A1(decode_regfile_fpregs_25__10_), .A2(n13317), .ZN(n2038)
         );
  NAND2_X2 U3645 ( .A1(decode_regfile_fpregs_25__0_), .A2(n13318), .ZN(n2039)
         );
  NAND2_X2 U3646 ( .A1(n1973), .A2(n800), .ZN(n2007) );
  NAND2_X2 U3648 ( .A1(decode_regfile_fpregs_24__9_), .A2(n13312), .ZN(n2041)
         );
  NAND2_X2 U3650 ( .A1(decode_regfile_fpregs_24__8_), .A2(n2040), .ZN(n2042)
         );
  NAND2_X2 U3652 ( .A1(decode_regfile_fpregs_24__7_), .A2(n2040), .ZN(n2043)
         );
  NAND2_X2 U3654 ( .A1(decode_regfile_fpregs_24__6_), .A2(n2040), .ZN(n2044)
         );
  NAND2_X2 U3656 ( .A1(decode_regfile_fpregs_24__5_), .A2(n2040), .ZN(n2045)
         );
  NAND2_X2 U3658 ( .A1(decode_regfile_fpregs_24__4_), .A2(n2040), .ZN(n2046)
         );
  NAND2_X2 U3660 ( .A1(decode_regfile_fpregs_24__3_), .A2(n2040), .ZN(n2047)
         );
  NAND2_X2 U3662 ( .A1(decode_regfile_fpregs_24__31_), .A2(n2040), .ZN(n2048)
         );
  NAND2_X2 U3664 ( .A1(decode_regfile_fpregs_24__30_), .A2(n13313), .ZN(n2049)
         );
  NAND2_X2 U3666 ( .A1(decode_regfile_fpregs_24__2_), .A2(n13313), .ZN(n2050)
         );
  NAND2_X2 U3668 ( .A1(decode_regfile_fpregs_24__29_), .A2(n13313), .ZN(n2051)
         );
  NAND2_X2 U3670 ( .A1(decode_regfile_fpregs_24__28_), .A2(n13313), .ZN(n2052)
         );
  NAND2_X2 U3672 ( .A1(decode_regfile_fpregs_24__27_), .A2(n13313), .ZN(n2053)
         );
  NAND2_X2 U3674 ( .A1(decode_regfile_fpregs_24__26_), .A2(n13313), .ZN(n2054)
         );
  NAND2_X2 U3676 ( .A1(decode_regfile_fpregs_24__25_), .A2(n13313), .ZN(n2055)
         );
  NAND2_X2 U3678 ( .A1(decode_regfile_fpregs_24__24_), .A2(n13313), .ZN(n2056)
         );
  NAND2_X2 U3680 ( .A1(decode_regfile_fpregs_24__23_), .A2(n13313), .ZN(n2057)
         );
  NAND2_X2 U3682 ( .A1(decode_regfile_fpregs_24__22_), .A2(n13313), .ZN(n2058)
         );
  NAND2_X2 U3684 ( .A1(decode_regfile_fpregs_24__21_), .A2(n13313), .ZN(n2059)
         );
  NAND2_X2 U3686 ( .A1(decode_regfile_fpregs_24__20_), .A2(n13313), .ZN(n2060)
         );
  NAND2_X2 U3688 ( .A1(decode_regfile_fpregs_24__1_), .A2(n13313), .ZN(n2061)
         );
  NAND2_X2 U3690 ( .A1(decode_regfile_fpregs_24__19_), .A2(n13313), .ZN(n2062)
         );
  NAND2_X2 U3692 ( .A1(decode_regfile_fpregs_24__18_), .A2(n13313), .ZN(n2063)
         );
  NAND2_X2 U3694 ( .A1(decode_regfile_fpregs_24__17_), .A2(n13313), .ZN(n2064)
         );
  NAND2_X2 U3696 ( .A1(decode_regfile_fpregs_24__16_), .A2(n13312), .ZN(n2065)
         );
  NAND2_X2 U3698 ( .A1(decode_regfile_fpregs_24__15_), .A2(n13312), .ZN(n2066)
         );
  NAND2_X2 U3700 ( .A1(decode_regfile_fpregs_24__14_), .A2(n13313), .ZN(n2067)
         );
  NAND2_X2 U3702 ( .A1(decode_regfile_fpregs_24__13_), .A2(n13312), .ZN(n2068)
         );
  NAND2_X2 U3704 ( .A1(decode_regfile_fpregs_24__12_), .A2(n13312), .ZN(n2069)
         );
  NAND2_X2 U3706 ( .A1(decode_regfile_fpregs_24__11_), .A2(n13313), .ZN(n2070)
         );
  NAND2_X2 U3708 ( .A1(decode_regfile_fpregs_24__10_), .A2(n13312), .ZN(n2071)
         );
  NAND2_X2 U3710 ( .A1(decode_regfile_fpregs_24__0_), .A2(n13313), .ZN(n2072)
         );
  NAND2_X2 U3711 ( .A1(n1973), .A2(n834), .ZN(n2040) );
  AND2_X2 U3712 ( .A1(n1939), .A2(n461), .ZN(n1973) );
  NAND2_X2 U3714 ( .A1(decode_regfile_fpregs_23__9_), .A2(n13307), .ZN(n2074)
         );
  NAND2_X2 U3716 ( .A1(decode_regfile_fpregs_23__8_), .A2(n13309), .ZN(n2075)
         );
  NAND2_X2 U3718 ( .A1(decode_regfile_fpregs_23__7_), .A2(n13309), .ZN(n2076)
         );
  NAND2_X2 U3720 ( .A1(decode_regfile_fpregs_23__6_), .A2(n13309), .ZN(n2077)
         );
  NAND2_X2 U3722 ( .A1(decode_regfile_fpregs_23__5_), .A2(n13309), .ZN(n2078)
         );
  NAND2_X2 U3724 ( .A1(decode_regfile_fpregs_23__4_), .A2(n13309), .ZN(n2079)
         );
  NAND2_X2 U3726 ( .A1(decode_regfile_fpregs_23__3_), .A2(n13309), .ZN(n2080)
         );
  NAND2_X2 U3728 ( .A1(decode_regfile_fpregs_23__31_), .A2(n13309), .ZN(n2081)
         );
  NAND2_X2 U3730 ( .A1(decode_regfile_fpregs_23__30_), .A2(n13308), .ZN(n2082)
         );
  NAND2_X2 U3732 ( .A1(decode_regfile_fpregs_23__2_), .A2(n13308), .ZN(n2083)
         );
  NAND2_X2 U3734 ( .A1(decode_regfile_fpregs_23__29_), .A2(n13308), .ZN(n2084)
         );
  NAND2_X2 U3736 ( .A1(decode_regfile_fpregs_23__28_), .A2(n13308), .ZN(n2085)
         );
  NAND2_X2 U3738 ( .A1(decode_regfile_fpregs_23__27_), .A2(n13308), .ZN(n2086)
         );
  NAND2_X2 U3740 ( .A1(decode_regfile_fpregs_23__26_), .A2(n13308), .ZN(n2087)
         );
  NAND2_X2 U3742 ( .A1(decode_regfile_fpregs_23__25_), .A2(n13308), .ZN(n2088)
         );
  NAND2_X2 U3744 ( .A1(decode_regfile_fpregs_23__24_), .A2(n13308), .ZN(n2089)
         );
  NAND2_X2 U3746 ( .A1(decode_regfile_fpregs_23__23_), .A2(n13308), .ZN(n2090)
         );
  NAND2_X2 U3748 ( .A1(decode_regfile_fpregs_23__22_), .A2(n13308), .ZN(n2091)
         );
  NAND2_X2 U3750 ( .A1(decode_regfile_fpregs_23__21_), .A2(n13308), .ZN(n2092)
         );
  NAND2_X2 U3752 ( .A1(decode_regfile_fpregs_23__20_), .A2(n13308), .ZN(n2093)
         );
  NAND2_X2 U3754 ( .A1(decode_regfile_fpregs_23__1_), .A2(n13308), .ZN(n2094)
         );
  NAND2_X2 U3756 ( .A1(decode_regfile_fpregs_23__19_), .A2(n13308), .ZN(n2095)
         );
  NAND2_X2 U3758 ( .A1(decode_regfile_fpregs_23__18_), .A2(n13308), .ZN(n2096)
         );
  NAND2_X2 U3760 ( .A1(decode_regfile_fpregs_23__17_), .A2(n13308), .ZN(n2097)
         );
  NAND2_X2 U3762 ( .A1(decode_regfile_fpregs_23__16_), .A2(n13307), .ZN(n2098)
         );
  NAND2_X2 U3764 ( .A1(decode_regfile_fpregs_23__15_), .A2(n13307), .ZN(n2099)
         );
  NAND2_X2 U3766 ( .A1(decode_regfile_fpregs_23__14_), .A2(n13308), .ZN(n2100)
         );
  NAND2_X2 U3768 ( .A1(decode_regfile_fpregs_23__13_), .A2(n13307), .ZN(n2101)
         );
  NAND2_X2 U3770 ( .A1(decode_regfile_fpregs_23__12_), .A2(n13307), .ZN(n2102)
         );
  NAND2_X2 U3772 ( .A1(decode_regfile_fpregs_23__11_), .A2(n13308), .ZN(n2103)
         );
  NAND2_X2 U3774 ( .A1(decode_regfile_fpregs_23__10_), .A2(n13307), .ZN(n2104)
         );
  NAND2_X2 U3776 ( .A1(decode_regfile_fpregs_23__0_), .A2(n13308), .ZN(n2105)
         );
  NAND2_X2 U3779 ( .A1(decode_regfile_fpregs_22__9_), .A2(n13302), .ZN(n2108)
         );
  NAND2_X2 U3781 ( .A1(decode_regfile_fpregs_22__8_), .A2(n13304), .ZN(n2109)
         );
  NAND2_X2 U3783 ( .A1(decode_regfile_fpregs_22__7_), .A2(n13304), .ZN(n2110)
         );
  NAND2_X2 U3785 ( .A1(decode_regfile_fpregs_22__6_), .A2(n13304), .ZN(n2111)
         );
  NAND2_X2 U3787 ( .A1(decode_regfile_fpregs_22__5_), .A2(n13304), .ZN(n2112)
         );
  NAND2_X2 U3789 ( .A1(decode_regfile_fpregs_22__4_), .A2(n13304), .ZN(n2113)
         );
  NAND2_X2 U3791 ( .A1(decode_regfile_fpregs_22__3_), .A2(n13304), .ZN(n2114)
         );
  NAND2_X2 U3793 ( .A1(decode_regfile_fpregs_22__31_), .A2(n13304), .ZN(n2115)
         );
  NAND2_X2 U3795 ( .A1(decode_regfile_fpregs_22__30_), .A2(n13303), .ZN(n2116)
         );
  NAND2_X2 U3797 ( .A1(decode_regfile_fpregs_22__2_), .A2(n13303), .ZN(n2117)
         );
  NAND2_X2 U3799 ( .A1(decode_regfile_fpregs_22__29_), .A2(n13303), .ZN(n2118)
         );
  NAND2_X2 U3801 ( .A1(decode_regfile_fpregs_22__28_), .A2(n13303), .ZN(n2119)
         );
  NAND2_X2 U3803 ( .A1(decode_regfile_fpregs_22__27_), .A2(n13303), .ZN(n2120)
         );
  NAND2_X2 U3805 ( .A1(decode_regfile_fpregs_22__26_), .A2(n13303), .ZN(n2121)
         );
  NAND2_X2 U3807 ( .A1(decode_regfile_fpregs_22__25_), .A2(n13303), .ZN(n2122)
         );
  NAND2_X2 U3809 ( .A1(decode_regfile_fpregs_22__24_), .A2(n13303), .ZN(n2123)
         );
  NAND2_X2 U3811 ( .A1(decode_regfile_fpregs_22__23_), .A2(n13303), .ZN(n2124)
         );
  NAND2_X2 U3813 ( .A1(decode_regfile_fpregs_22__22_), .A2(n13303), .ZN(n2125)
         );
  NAND2_X2 U3815 ( .A1(decode_regfile_fpregs_22__21_), .A2(n13303), .ZN(n2126)
         );
  NAND2_X2 U3817 ( .A1(decode_regfile_fpregs_22__20_), .A2(n13303), .ZN(n2127)
         );
  NAND2_X2 U3819 ( .A1(decode_regfile_fpregs_22__1_), .A2(n13303), .ZN(n2128)
         );
  NAND2_X2 U3821 ( .A1(decode_regfile_fpregs_22__19_), .A2(n13303), .ZN(n2129)
         );
  NAND2_X2 U3823 ( .A1(decode_regfile_fpregs_22__18_), .A2(n13303), .ZN(n2130)
         );
  NAND2_X2 U3825 ( .A1(decode_regfile_fpregs_22__17_), .A2(n13303), .ZN(n2131)
         );
  NAND2_X2 U3827 ( .A1(decode_regfile_fpregs_22__16_), .A2(n13302), .ZN(n2132)
         );
  NAND2_X2 U3829 ( .A1(decode_regfile_fpregs_22__15_), .A2(n13302), .ZN(n2133)
         );
  NAND2_X2 U3831 ( .A1(decode_regfile_fpregs_22__14_), .A2(n13303), .ZN(n2134)
         );
  NAND2_X2 U3833 ( .A1(decode_regfile_fpregs_22__13_), .A2(n13302), .ZN(n2135)
         );
  NAND2_X2 U3835 ( .A1(decode_regfile_fpregs_22__12_), .A2(n13302), .ZN(n2136)
         );
  NAND2_X2 U3837 ( .A1(decode_regfile_fpregs_22__11_), .A2(n13303), .ZN(n2137)
         );
  NAND2_X2 U3839 ( .A1(decode_regfile_fpregs_22__10_), .A2(n13302), .ZN(n2138)
         );
  NAND2_X2 U3841 ( .A1(decode_regfile_fpregs_22__0_), .A2(n13303), .ZN(n2139)
         );
  NAND2_X2 U3844 ( .A1(decode_regfile_fpregs_21__9_), .A2(n13297), .ZN(n2141)
         );
  NAND2_X2 U3846 ( .A1(decode_regfile_fpregs_21__8_), .A2(n2140), .ZN(n2142)
         );
  NAND2_X2 U3848 ( .A1(decode_regfile_fpregs_21__7_), .A2(n2140), .ZN(n2143)
         );
  NAND2_X2 U3850 ( .A1(decode_regfile_fpregs_21__6_), .A2(n2140), .ZN(n2144)
         );
  NAND2_X2 U3852 ( .A1(decode_regfile_fpregs_21__5_), .A2(n2140), .ZN(n2145)
         );
  NAND2_X2 U3854 ( .A1(decode_regfile_fpregs_21__4_), .A2(n2140), .ZN(n2146)
         );
  NAND2_X2 U3856 ( .A1(decode_regfile_fpregs_21__3_), .A2(n2140), .ZN(n2147)
         );
  NAND2_X2 U3858 ( .A1(decode_regfile_fpregs_21__31_), .A2(n2140), .ZN(n2148)
         );
  NAND2_X2 U3860 ( .A1(decode_regfile_fpregs_21__30_), .A2(n13298), .ZN(n2149)
         );
  NAND2_X2 U3862 ( .A1(decode_regfile_fpregs_21__2_), .A2(n13298), .ZN(n2150)
         );
  NAND2_X2 U3864 ( .A1(decode_regfile_fpregs_21__29_), .A2(n13298), .ZN(n2151)
         );
  NAND2_X2 U3866 ( .A1(decode_regfile_fpregs_21__28_), .A2(n13298), .ZN(n2152)
         );
  NAND2_X2 U3868 ( .A1(decode_regfile_fpregs_21__27_), .A2(n13298), .ZN(n2153)
         );
  NAND2_X2 U3870 ( .A1(decode_regfile_fpregs_21__26_), .A2(n13298), .ZN(n2154)
         );
  NAND2_X2 U3872 ( .A1(decode_regfile_fpregs_21__25_), .A2(n13298), .ZN(n2155)
         );
  NAND2_X2 U3874 ( .A1(decode_regfile_fpregs_21__24_), .A2(n13298), .ZN(n2156)
         );
  NAND2_X2 U3876 ( .A1(decode_regfile_fpregs_21__23_), .A2(n13298), .ZN(n2157)
         );
  NAND2_X2 U3878 ( .A1(decode_regfile_fpregs_21__22_), .A2(n13298), .ZN(n2158)
         );
  NAND2_X2 U3880 ( .A1(decode_regfile_fpregs_21__21_), .A2(n13298), .ZN(n2159)
         );
  NAND2_X2 U3882 ( .A1(decode_regfile_fpregs_21__20_), .A2(n13298), .ZN(n2160)
         );
  NAND2_X2 U3884 ( .A1(decode_regfile_fpregs_21__1_), .A2(n13298), .ZN(n2161)
         );
  NAND2_X2 U3886 ( .A1(decode_regfile_fpregs_21__19_), .A2(n13298), .ZN(n2162)
         );
  NAND2_X2 U3888 ( .A1(decode_regfile_fpregs_21__18_), .A2(n13298), .ZN(n2163)
         );
  NAND2_X2 U3890 ( .A1(decode_regfile_fpregs_21__17_), .A2(n13298), .ZN(n2164)
         );
  NAND2_X2 U3892 ( .A1(decode_regfile_fpregs_21__16_), .A2(n13297), .ZN(n2165)
         );
  NAND2_X2 U3894 ( .A1(decode_regfile_fpregs_21__15_), .A2(n13297), .ZN(n2166)
         );
  NAND2_X2 U3896 ( .A1(decode_regfile_fpregs_21__14_), .A2(n13298), .ZN(n2167)
         );
  NAND2_X2 U3898 ( .A1(decode_regfile_fpregs_21__13_), .A2(n13297), .ZN(n2168)
         );
  NAND2_X2 U3900 ( .A1(decode_regfile_fpregs_21__12_), .A2(n13297), .ZN(n2169)
         );
  NAND2_X2 U3902 ( .A1(decode_regfile_fpregs_21__11_), .A2(n13298), .ZN(n2170)
         );
  NAND2_X2 U3904 ( .A1(decode_regfile_fpregs_21__10_), .A2(n13297), .ZN(n2171)
         );
  NAND2_X2 U3906 ( .A1(decode_regfile_fpregs_21__0_), .A2(n13298), .ZN(n2172)
         );
  NAND2_X2 U3907 ( .A1(n2106), .A2(n800), .ZN(n2140) );
  NAND2_X2 U3909 ( .A1(decode_regfile_fpregs_20__9_), .A2(n13292), .ZN(n2174)
         );
  NAND2_X2 U3911 ( .A1(decode_regfile_fpregs_20__8_), .A2(n2173), .ZN(n2175)
         );
  NAND2_X2 U3913 ( .A1(decode_regfile_fpregs_20__7_), .A2(n2173), .ZN(n2176)
         );
  NAND2_X2 U3915 ( .A1(decode_regfile_fpregs_20__6_), .A2(n2173), .ZN(n2177)
         );
  NAND2_X2 U3917 ( .A1(decode_regfile_fpregs_20__5_), .A2(n2173), .ZN(n2178)
         );
  NAND2_X2 U3919 ( .A1(decode_regfile_fpregs_20__4_), .A2(n2173), .ZN(n2179)
         );
  NAND2_X2 U3921 ( .A1(decode_regfile_fpregs_20__3_), .A2(n2173), .ZN(n2180)
         );
  NAND2_X2 U3923 ( .A1(decode_regfile_fpregs_20__31_), .A2(n2173), .ZN(n2181)
         );
  NAND2_X2 U3925 ( .A1(decode_regfile_fpregs_20__30_), .A2(n13293), .ZN(n2182)
         );
  NAND2_X2 U3927 ( .A1(decode_regfile_fpregs_20__2_), .A2(n13293), .ZN(n2183)
         );
  NAND2_X2 U3929 ( .A1(decode_regfile_fpregs_20__29_), .A2(n13293), .ZN(n2184)
         );
  NAND2_X2 U3931 ( .A1(decode_regfile_fpregs_20__28_), .A2(n13293), .ZN(n2185)
         );
  NAND2_X2 U3933 ( .A1(decode_regfile_fpregs_20__27_), .A2(n13293), .ZN(n2186)
         );
  NAND2_X2 U3935 ( .A1(decode_regfile_fpregs_20__26_), .A2(n13293), .ZN(n2187)
         );
  NAND2_X2 U3937 ( .A1(decode_regfile_fpregs_20__25_), .A2(n13293), .ZN(n2188)
         );
  NAND2_X2 U3939 ( .A1(decode_regfile_fpregs_20__24_), .A2(n13293), .ZN(n2189)
         );
  NAND2_X2 U3941 ( .A1(decode_regfile_fpregs_20__23_), .A2(n13293), .ZN(n2190)
         );
  NAND2_X2 U3943 ( .A1(decode_regfile_fpregs_20__22_), .A2(n13293), .ZN(n2191)
         );
  NAND2_X2 U3945 ( .A1(decode_regfile_fpregs_20__21_), .A2(n13293), .ZN(n2192)
         );
  NAND2_X2 U3947 ( .A1(decode_regfile_fpregs_20__20_), .A2(n13293), .ZN(n2193)
         );
  NAND2_X2 U3949 ( .A1(decode_regfile_fpregs_20__1_), .A2(n13293), .ZN(n2194)
         );
  NAND2_X2 U3951 ( .A1(decode_regfile_fpregs_20__19_), .A2(n13293), .ZN(n2195)
         );
  NAND2_X2 U3953 ( .A1(decode_regfile_fpregs_20__18_), .A2(n13293), .ZN(n2196)
         );
  NAND2_X2 U3955 ( .A1(decode_regfile_fpregs_20__17_), .A2(n13293), .ZN(n2197)
         );
  NAND2_X2 U3957 ( .A1(decode_regfile_fpregs_20__16_), .A2(n13292), .ZN(n2198)
         );
  NAND2_X2 U3959 ( .A1(decode_regfile_fpregs_20__15_), .A2(n13292), .ZN(n2199)
         );
  NAND2_X2 U3961 ( .A1(decode_regfile_fpregs_20__14_), .A2(n13293), .ZN(n2200)
         );
  NAND2_X2 U3963 ( .A1(decode_regfile_fpregs_20__13_), .A2(n13292), .ZN(n2201)
         );
  NAND2_X2 U3965 ( .A1(decode_regfile_fpregs_20__12_), .A2(n13292), .ZN(n2202)
         );
  NAND2_X2 U3967 ( .A1(decode_regfile_fpregs_20__11_), .A2(n13293), .ZN(n2203)
         );
  NAND2_X2 U3969 ( .A1(decode_regfile_fpregs_20__10_), .A2(n13292), .ZN(n2204)
         );
  NAND2_X2 U3971 ( .A1(decode_regfile_fpregs_20__0_), .A2(n13293), .ZN(n2205)
         );
  NAND2_X2 U3972 ( .A1(n2106), .A2(n834), .ZN(n2173) );
  AND2_X2 U3973 ( .A1(n1939), .A2(n530), .ZN(n2106) );
  NAND2_X2 U3976 ( .A1(decode_regfile_fpregs_1__9_), .A2(n13287), .ZN(n2208)
         );
  NAND2_X2 U3978 ( .A1(decode_regfile_fpregs_1__8_), .A2(n2207), .ZN(n2209) );
  NAND2_X2 U3980 ( .A1(decode_regfile_fpregs_1__7_), .A2(n2207), .ZN(n2210) );
  NAND2_X2 U3982 ( .A1(decode_regfile_fpregs_1__6_), .A2(n2207), .ZN(n2211) );
  NAND2_X2 U3984 ( .A1(decode_regfile_fpregs_1__5_), .A2(n2207), .ZN(n2212) );
  NAND2_X2 U3986 ( .A1(decode_regfile_fpregs_1__4_), .A2(n2207), .ZN(n2213) );
  NAND2_X2 U3988 ( .A1(decode_regfile_fpregs_1__3_), .A2(n2207), .ZN(n2214) );
  NAND2_X2 U3990 ( .A1(decode_regfile_fpregs_1__31_), .A2(n2207), .ZN(n2215)
         );
  NAND2_X2 U3992 ( .A1(decode_regfile_fpregs_1__30_), .A2(n13288), .ZN(n2216)
         );
  NAND2_X2 U3994 ( .A1(decode_regfile_fpregs_1__2_), .A2(n13288), .ZN(n2217)
         );
  NAND2_X2 U3996 ( .A1(decode_regfile_fpregs_1__29_), .A2(n13288), .ZN(n2218)
         );
  NAND2_X2 U3998 ( .A1(decode_regfile_fpregs_1__28_), .A2(n13288), .ZN(n2219)
         );
  NAND2_X2 U4000 ( .A1(decode_regfile_fpregs_1__27_), .A2(n13288), .ZN(n2220)
         );
  NAND2_X2 U4002 ( .A1(decode_regfile_fpregs_1__26_), .A2(n13288), .ZN(n2221)
         );
  NAND2_X2 U4004 ( .A1(decode_regfile_fpregs_1__25_), .A2(n13288), .ZN(n2222)
         );
  NAND2_X2 U4006 ( .A1(decode_regfile_fpregs_1__24_), .A2(n13288), .ZN(n2223)
         );
  NAND2_X2 U4008 ( .A1(decode_regfile_fpregs_1__23_), .A2(n13288), .ZN(n2224)
         );
  NAND2_X2 U4010 ( .A1(decode_regfile_fpregs_1__22_), .A2(n13288), .ZN(n2225)
         );
  NAND2_X2 U4012 ( .A1(decode_regfile_fpregs_1__21_), .A2(n13288), .ZN(n2226)
         );
  NAND2_X2 U4014 ( .A1(decode_regfile_fpregs_1__20_), .A2(n13288), .ZN(n2227)
         );
  NAND2_X2 U4016 ( .A1(decode_regfile_fpregs_1__1_), .A2(n13288), .ZN(n2228)
         );
  NAND2_X2 U4018 ( .A1(decode_regfile_fpregs_1__19_), .A2(n13288), .ZN(n2229)
         );
  NAND2_X2 U4020 ( .A1(decode_regfile_fpregs_1__18_), .A2(n13288), .ZN(n2230)
         );
  NAND2_X2 U4022 ( .A1(decode_regfile_fpregs_1__17_), .A2(n13288), .ZN(n2231)
         );
  NAND2_X2 U4024 ( .A1(decode_regfile_fpregs_1__16_), .A2(n13287), .ZN(n2232)
         );
  NAND2_X2 U4026 ( .A1(decode_regfile_fpregs_1__15_), .A2(n13287), .ZN(n2233)
         );
  NAND2_X2 U4028 ( .A1(decode_regfile_fpregs_1__14_), .A2(n13288), .ZN(n2234)
         );
  NAND2_X2 U4030 ( .A1(decode_regfile_fpregs_1__13_), .A2(n13287), .ZN(n2235)
         );
  NAND2_X2 U4032 ( .A1(decode_regfile_fpregs_1__12_), .A2(n13287), .ZN(n2236)
         );
  NAND2_X2 U4034 ( .A1(decode_regfile_fpregs_1__11_), .A2(n13288), .ZN(n2237)
         );
  NAND2_X2 U4036 ( .A1(decode_regfile_fpregs_1__10_), .A2(n13287), .ZN(n2238)
         );
  NAND2_X2 U4038 ( .A1(decode_regfile_fpregs_1__0_), .A2(n13288), .ZN(n2239)
         );
  NAND2_X2 U4039 ( .A1(n1772), .A2(n800), .ZN(n2207) );
  NAND2_X2 U4041 ( .A1(decode_regfile_fpregs_19__9_), .A2(n13282), .ZN(n2241)
         );
  NAND2_X2 U4043 ( .A1(decode_regfile_fpregs_19__8_), .A2(n13284), .ZN(n2242)
         );
  NAND2_X2 U4045 ( .A1(decode_regfile_fpregs_19__7_), .A2(n13284), .ZN(n2243)
         );
  NAND2_X2 U4047 ( .A1(decode_regfile_fpregs_19__6_), .A2(n13284), .ZN(n2244)
         );
  NAND2_X2 U4049 ( .A1(decode_regfile_fpregs_19__5_), .A2(n13284), .ZN(n2245)
         );
  NAND2_X2 U4051 ( .A1(decode_regfile_fpregs_19__4_), .A2(n13284), .ZN(n2246)
         );
  NAND2_X2 U4053 ( .A1(decode_regfile_fpregs_19__3_), .A2(n13284), .ZN(n2247)
         );
  NAND2_X2 U4055 ( .A1(decode_regfile_fpregs_19__31_), .A2(n13284), .ZN(n2248)
         );
  NAND2_X2 U4057 ( .A1(decode_regfile_fpregs_19__30_), .A2(n13283), .ZN(n2249)
         );
  NAND2_X2 U4059 ( .A1(decode_regfile_fpregs_19__2_), .A2(n13283), .ZN(n2250)
         );
  NAND2_X2 U4061 ( .A1(decode_regfile_fpregs_19__29_), .A2(n13283), .ZN(n2251)
         );
  NAND2_X2 U4063 ( .A1(decode_regfile_fpregs_19__28_), .A2(n13283), .ZN(n2252)
         );
  NAND2_X2 U4065 ( .A1(decode_regfile_fpregs_19__27_), .A2(n13283), .ZN(n2253)
         );
  NAND2_X2 U4067 ( .A1(decode_regfile_fpregs_19__26_), .A2(n13283), .ZN(n2254)
         );
  NAND2_X2 U4069 ( .A1(decode_regfile_fpregs_19__25_), .A2(n13283), .ZN(n2255)
         );
  NAND2_X2 U4071 ( .A1(decode_regfile_fpregs_19__24_), .A2(n13283), .ZN(n2256)
         );
  NAND2_X2 U4073 ( .A1(decode_regfile_fpregs_19__23_), .A2(n13283), .ZN(n2257)
         );
  NAND2_X2 U4075 ( .A1(decode_regfile_fpregs_19__22_), .A2(n13283), .ZN(n2258)
         );
  NAND2_X2 U4077 ( .A1(decode_regfile_fpregs_19__21_), .A2(n13283), .ZN(n2259)
         );
  NAND2_X2 U4079 ( .A1(decode_regfile_fpregs_19__20_), .A2(n13283), .ZN(n2260)
         );
  NAND2_X2 U4081 ( .A1(decode_regfile_fpregs_19__1_), .A2(n13283), .ZN(n2261)
         );
  NAND2_X2 U4083 ( .A1(decode_regfile_fpregs_19__19_), .A2(n13283), .ZN(n2262)
         );
  NAND2_X2 U4085 ( .A1(decode_regfile_fpregs_19__18_), .A2(n13283), .ZN(n2263)
         );
  NAND2_X2 U4087 ( .A1(decode_regfile_fpregs_19__17_), .A2(n13283), .ZN(n2264)
         );
  NAND2_X2 U4089 ( .A1(decode_regfile_fpregs_19__16_), .A2(n13282), .ZN(n2265)
         );
  NAND2_X2 U4091 ( .A1(decode_regfile_fpregs_19__15_), .A2(n13282), .ZN(n2266)
         );
  NAND2_X2 U4093 ( .A1(decode_regfile_fpregs_19__14_), .A2(n13283), .ZN(n2267)
         );
  NAND2_X2 U4095 ( .A1(decode_regfile_fpregs_19__13_), .A2(n13282), .ZN(n2268)
         );
  NAND2_X2 U4097 ( .A1(decode_regfile_fpregs_19__12_), .A2(n13282), .ZN(n2269)
         );
  NAND2_X2 U4099 ( .A1(decode_regfile_fpregs_19__11_), .A2(n13283), .ZN(n2270)
         );
  NAND2_X2 U4101 ( .A1(decode_regfile_fpregs_19__10_), .A2(n13282), .ZN(n2271)
         );
  NAND2_X2 U4103 ( .A1(decode_regfile_fpregs_19__0_), .A2(n13283), .ZN(n2272)
         );
  NAND2_X2 U4106 ( .A1(decode_regfile_fpregs_18__9_), .A2(n13277), .ZN(n2275)
         );
  NAND2_X2 U4108 ( .A1(decode_regfile_fpregs_18__8_), .A2(n13279), .ZN(n2276)
         );
  NAND2_X2 U4110 ( .A1(decode_regfile_fpregs_18__7_), .A2(n13279), .ZN(n2277)
         );
  NAND2_X2 U4112 ( .A1(decode_regfile_fpregs_18__6_), .A2(n13279), .ZN(n2278)
         );
  NAND2_X2 U4114 ( .A1(decode_regfile_fpregs_18__5_), .A2(n13279), .ZN(n2279)
         );
  NAND2_X2 U4116 ( .A1(decode_regfile_fpregs_18__4_), .A2(n13279), .ZN(n2280)
         );
  NAND2_X2 U4118 ( .A1(decode_regfile_fpregs_18__3_), .A2(n13279), .ZN(n2281)
         );
  NAND2_X2 U4120 ( .A1(decode_regfile_fpregs_18__31_), .A2(n13279), .ZN(n2282)
         );
  NAND2_X2 U4122 ( .A1(decode_regfile_fpregs_18__30_), .A2(n13278), .ZN(n2283)
         );
  NAND2_X2 U4124 ( .A1(decode_regfile_fpregs_18__2_), .A2(n13278), .ZN(n2284)
         );
  NAND2_X2 U4126 ( .A1(decode_regfile_fpregs_18__29_), .A2(n13278), .ZN(n2285)
         );
  NAND2_X2 U4128 ( .A1(decode_regfile_fpregs_18__28_), .A2(n13278), .ZN(n2286)
         );
  NAND2_X2 U4130 ( .A1(decode_regfile_fpregs_18__27_), .A2(n13278), .ZN(n2287)
         );
  NAND2_X2 U4132 ( .A1(decode_regfile_fpregs_18__26_), .A2(n13278), .ZN(n2288)
         );
  NAND2_X2 U4134 ( .A1(decode_regfile_fpregs_18__25_), .A2(n13278), .ZN(n2289)
         );
  NAND2_X2 U4136 ( .A1(decode_regfile_fpregs_18__24_), .A2(n13278), .ZN(n2290)
         );
  NAND2_X2 U4138 ( .A1(decode_regfile_fpregs_18__23_), .A2(n13278), .ZN(n2291)
         );
  NAND2_X2 U4140 ( .A1(decode_regfile_fpregs_18__22_), .A2(n13278), .ZN(n2292)
         );
  NAND2_X2 U4142 ( .A1(decode_regfile_fpregs_18__21_), .A2(n13278), .ZN(n2293)
         );
  NAND2_X2 U4144 ( .A1(decode_regfile_fpregs_18__20_), .A2(n13278), .ZN(n2294)
         );
  NAND2_X2 U4146 ( .A1(decode_regfile_fpregs_18__1_), .A2(n13278), .ZN(n2295)
         );
  NAND2_X2 U4148 ( .A1(decode_regfile_fpregs_18__19_), .A2(n13278), .ZN(n2296)
         );
  NAND2_X2 U4150 ( .A1(decode_regfile_fpregs_18__18_), .A2(n13278), .ZN(n2297)
         );
  NAND2_X2 U4152 ( .A1(decode_regfile_fpregs_18__17_), .A2(n13278), .ZN(n2298)
         );
  NAND2_X2 U4154 ( .A1(decode_regfile_fpregs_18__16_), .A2(n13277), .ZN(n2299)
         );
  NAND2_X2 U4156 ( .A1(decode_regfile_fpregs_18__15_), .A2(n13277), .ZN(n2300)
         );
  NAND2_X2 U4158 ( .A1(decode_regfile_fpregs_18__14_), .A2(n13278), .ZN(n2301)
         );
  NAND2_X2 U4160 ( .A1(decode_regfile_fpregs_18__13_), .A2(n13277), .ZN(n2302)
         );
  NAND2_X2 U4162 ( .A1(decode_regfile_fpregs_18__12_), .A2(n13277), .ZN(n2303)
         );
  NAND2_X2 U4164 ( .A1(decode_regfile_fpregs_18__11_), .A2(n13278), .ZN(n2304)
         );
  NAND2_X2 U4166 ( .A1(decode_regfile_fpregs_18__10_), .A2(n13277), .ZN(n2305)
         );
  NAND2_X2 U4168 ( .A1(decode_regfile_fpregs_18__0_), .A2(n13278), .ZN(n2306)
         );
  NAND2_X2 U4171 ( .A1(decode_regfile_fpregs_17__9_), .A2(n13272), .ZN(n2308)
         );
  NAND2_X2 U4173 ( .A1(decode_regfile_fpregs_17__8_), .A2(n2307), .ZN(n2309)
         );
  NAND2_X2 U4175 ( .A1(decode_regfile_fpregs_17__7_), .A2(n2307), .ZN(n2310)
         );
  NAND2_X2 U4177 ( .A1(decode_regfile_fpregs_17__6_), .A2(n2307), .ZN(n2311)
         );
  NAND2_X2 U4179 ( .A1(decode_regfile_fpregs_17__5_), .A2(n2307), .ZN(n2312)
         );
  NAND2_X2 U4181 ( .A1(decode_regfile_fpregs_17__4_), .A2(n2307), .ZN(n2313)
         );
  NAND2_X2 U4183 ( .A1(decode_regfile_fpregs_17__3_), .A2(n2307), .ZN(n2314)
         );
  NAND2_X2 U4185 ( .A1(decode_regfile_fpregs_17__31_), .A2(n2307), .ZN(n2315)
         );
  NAND2_X2 U4187 ( .A1(decode_regfile_fpregs_17__30_), .A2(n13273), .ZN(n2316)
         );
  NAND2_X2 U4189 ( .A1(decode_regfile_fpregs_17__2_), .A2(n13273), .ZN(n2317)
         );
  NAND2_X2 U4191 ( .A1(decode_regfile_fpregs_17__29_), .A2(n13273), .ZN(n2318)
         );
  NAND2_X2 U4193 ( .A1(decode_regfile_fpregs_17__28_), .A2(n13273), .ZN(n2319)
         );
  NAND2_X2 U4195 ( .A1(decode_regfile_fpregs_17__27_), .A2(n13273), .ZN(n2320)
         );
  NAND2_X2 U4197 ( .A1(decode_regfile_fpregs_17__26_), .A2(n13273), .ZN(n2321)
         );
  NAND2_X2 U4199 ( .A1(decode_regfile_fpregs_17__25_), .A2(n13273), .ZN(n2322)
         );
  NAND2_X2 U4201 ( .A1(decode_regfile_fpregs_17__24_), .A2(n13273), .ZN(n2323)
         );
  NAND2_X2 U4203 ( .A1(decode_regfile_fpregs_17__23_), .A2(n13273), .ZN(n2324)
         );
  NAND2_X2 U4205 ( .A1(decode_regfile_fpregs_17__22_), .A2(n13273), .ZN(n2325)
         );
  NAND2_X2 U4207 ( .A1(decode_regfile_fpregs_17__21_), .A2(n13273), .ZN(n2326)
         );
  NAND2_X2 U4209 ( .A1(decode_regfile_fpregs_17__20_), .A2(n13273), .ZN(n2327)
         );
  NAND2_X2 U4211 ( .A1(decode_regfile_fpregs_17__1_), .A2(n13273), .ZN(n2328)
         );
  NAND2_X2 U4213 ( .A1(decode_regfile_fpregs_17__19_), .A2(n13273), .ZN(n2329)
         );
  NAND2_X2 U4215 ( .A1(decode_regfile_fpregs_17__18_), .A2(n13273), .ZN(n2330)
         );
  NAND2_X2 U4217 ( .A1(decode_regfile_fpregs_17__17_), .A2(n13273), .ZN(n2331)
         );
  NAND2_X2 U4219 ( .A1(decode_regfile_fpregs_17__16_), .A2(n13272), .ZN(n2332)
         );
  NAND2_X2 U4221 ( .A1(decode_regfile_fpregs_17__15_), .A2(n13272), .ZN(n2333)
         );
  NAND2_X2 U4223 ( .A1(decode_regfile_fpregs_17__14_), .A2(n13273), .ZN(n2334)
         );
  NAND2_X2 U4225 ( .A1(decode_regfile_fpregs_17__13_), .A2(n13272), .ZN(n2335)
         );
  NAND2_X2 U4227 ( .A1(decode_regfile_fpregs_17__12_), .A2(n13272), .ZN(n2336)
         );
  NAND2_X2 U4229 ( .A1(decode_regfile_fpregs_17__11_), .A2(n13273), .ZN(n2337)
         );
  NAND2_X2 U4231 ( .A1(decode_regfile_fpregs_17__10_), .A2(n13272), .ZN(n2338)
         );
  NAND2_X2 U4233 ( .A1(decode_regfile_fpregs_17__0_), .A2(n13273), .ZN(n2339)
         );
  NAND2_X2 U4234 ( .A1(n2273), .A2(n800), .ZN(n2307) );
  NAND2_X2 U4236 ( .A1(decode_regfile_fpregs_16__9_), .A2(n13267), .ZN(n2341)
         );
  NAND2_X2 U4238 ( .A1(decode_regfile_fpregs_16__8_), .A2(n2340), .ZN(n2342)
         );
  NAND2_X2 U4240 ( .A1(decode_regfile_fpregs_16__7_), .A2(n2340), .ZN(n2343)
         );
  NAND2_X2 U4242 ( .A1(decode_regfile_fpregs_16__6_), .A2(n2340), .ZN(n2344)
         );
  NAND2_X2 U4244 ( .A1(decode_regfile_fpregs_16__5_), .A2(n2340), .ZN(n2345)
         );
  NAND2_X2 U4246 ( .A1(decode_regfile_fpregs_16__4_), .A2(n2340), .ZN(n2346)
         );
  NAND2_X2 U4248 ( .A1(decode_regfile_fpregs_16__3_), .A2(n2340), .ZN(n2347)
         );
  NAND2_X2 U4250 ( .A1(decode_regfile_fpregs_16__31_), .A2(n2340), .ZN(n2348)
         );
  NAND2_X2 U4252 ( .A1(decode_regfile_fpregs_16__30_), .A2(n13268), .ZN(n2349)
         );
  NAND2_X2 U4254 ( .A1(decode_regfile_fpregs_16__2_), .A2(n13268), .ZN(n2350)
         );
  NAND2_X2 U4256 ( .A1(decode_regfile_fpregs_16__29_), .A2(n13268), .ZN(n2351)
         );
  NAND2_X2 U4258 ( .A1(decode_regfile_fpregs_16__28_), .A2(n13268), .ZN(n2352)
         );
  NAND2_X2 U4260 ( .A1(decode_regfile_fpregs_16__27_), .A2(n13268), .ZN(n2353)
         );
  NAND2_X2 U4262 ( .A1(decode_regfile_fpregs_16__26_), .A2(n13268), .ZN(n2354)
         );
  NAND2_X2 U4264 ( .A1(decode_regfile_fpregs_16__25_), .A2(n13268), .ZN(n2355)
         );
  NAND2_X2 U4266 ( .A1(decode_regfile_fpregs_16__24_), .A2(n13268), .ZN(n2356)
         );
  NAND2_X2 U4268 ( .A1(decode_regfile_fpregs_16__23_), .A2(n13268), .ZN(n2357)
         );
  NAND2_X2 U4270 ( .A1(decode_regfile_fpregs_16__22_), .A2(n13268), .ZN(n2358)
         );
  NAND2_X2 U4272 ( .A1(decode_regfile_fpregs_16__21_), .A2(n13268), .ZN(n2359)
         );
  NAND2_X2 U4274 ( .A1(decode_regfile_fpregs_16__20_), .A2(n13268), .ZN(n2360)
         );
  NAND2_X2 U4276 ( .A1(decode_regfile_fpregs_16__1_), .A2(n13268), .ZN(n2361)
         );
  NAND2_X2 U4278 ( .A1(decode_regfile_fpregs_16__19_), .A2(n13268), .ZN(n2362)
         );
  NAND2_X2 U4280 ( .A1(decode_regfile_fpregs_16__18_), .A2(n13268), .ZN(n2363)
         );
  NAND2_X2 U4282 ( .A1(decode_regfile_fpregs_16__17_), .A2(n13268), .ZN(n2364)
         );
  NAND2_X2 U4284 ( .A1(decode_regfile_fpregs_16__16_), .A2(n13267), .ZN(n2365)
         );
  NAND2_X2 U4286 ( .A1(decode_regfile_fpregs_16__15_), .A2(n13267), .ZN(n2366)
         );
  NAND2_X2 U4288 ( .A1(decode_regfile_fpregs_16__14_), .A2(n13268), .ZN(n2367)
         );
  NAND2_X2 U4290 ( .A1(decode_regfile_fpregs_16__13_), .A2(n13267), .ZN(n2368)
         );
  NAND2_X2 U4292 ( .A1(decode_regfile_fpregs_16__12_), .A2(n13267), .ZN(n2369)
         );
  NAND2_X2 U4294 ( .A1(decode_regfile_fpregs_16__11_), .A2(n13268), .ZN(n2370)
         );
  NAND2_X2 U4296 ( .A1(decode_regfile_fpregs_16__10_), .A2(n13267), .ZN(n2371)
         );
  NAND2_X2 U4298 ( .A1(decode_regfile_fpregs_16__0_), .A2(n13268), .ZN(n2372)
         );
  NAND2_X2 U4299 ( .A1(n2273), .A2(n834), .ZN(n2340) );
  AND2_X2 U4300 ( .A1(n1939), .A2(n664), .ZN(n2273) );
  NAND2_X2 U4304 ( .A1(decode_regfile_fpregs_15__9_), .A2(n13262), .ZN(n2375)
         );
  NAND2_X2 U4306 ( .A1(decode_regfile_fpregs_15__8_), .A2(n13264), .ZN(n2376)
         );
  NAND2_X2 U4308 ( .A1(decode_regfile_fpregs_15__7_), .A2(n13264), .ZN(n2377)
         );
  NAND2_X2 U4310 ( .A1(decode_regfile_fpregs_15__6_), .A2(n13264), .ZN(n2378)
         );
  NAND2_X2 U4312 ( .A1(decode_regfile_fpregs_15__5_), .A2(n13264), .ZN(n2379)
         );
  NAND2_X2 U4314 ( .A1(decode_regfile_fpregs_15__4_), .A2(n13264), .ZN(n2380)
         );
  NAND2_X2 U4316 ( .A1(decode_regfile_fpregs_15__3_), .A2(n13264), .ZN(n2381)
         );
  NAND2_X2 U4318 ( .A1(decode_regfile_fpregs_15__31_), .A2(n13264), .ZN(n2382)
         );
  NAND2_X2 U4320 ( .A1(decode_regfile_fpregs_15__30_), .A2(n13263), .ZN(n2383)
         );
  NAND2_X2 U4322 ( .A1(decode_regfile_fpregs_15__2_), .A2(n13263), .ZN(n2384)
         );
  NAND2_X2 U4324 ( .A1(decode_regfile_fpregs_15__29_), .A2(n13263), .ZN(n2385)
         );
  NAND2_X2 U4326 ( .A1(decode_regfile_fpregs_15__28_), .A2(n13263), .ZN(n2386)
         );
  NAND2_X2 U4328 ( .A1(decode_regfile_fpregs_15__27_), .A2(n13263), .ZN(n2387)
         );
  NAND2_X2 U4330 ( .A1(decode_regfile_fpregs_15__26_), .A2(n13263), .ZN(n2388)
         );
  NAND2_X2 U4332 ( .A1(decode_regfile_fpregs_15__25_), .A2(n13263), .ZN(n2389)
         );
  NAND2_X2 U4334 ( .A1(decode_regfile_fpregs_15__24_), .A2(n13263), .ZN(n2390)
         );
  NAND2_X2 U4336 ( .A1(decode_regfile_fpregs_15__23_), .A2(n13263), .ZN(n2391)
         );
  NAND2_X2 U4338 ( .A1(decode_regfile_fpregs_15__22_), .A2(n13263), .ZN(n2392)
         );
  NAND2_X2 U4340 ( .A1(decode_regfile_fpregs_15__21_), .A2(n13263), .ZN(n2393)
         );
  NAND2_X2 U4342 ( .A1(decode_regfile_fpregs_15__20_), .A2(n13263), .ZN(n2394)
         );
  NAND2_X2 U4344 ( .A1(decode_regfile_fpregs_15__1_), .A2(n13263), .ZN(n2395)
         );
  NAND2_X2 U4346 ( .A1(decode_regfile_fpregs_15__19_), .A2(n13263), .ZN(n2396)
         );
  NAND2_X2 U4348 ( .A1(decode_regfile_fpregs_15__18_), .A2(n13263), .ZN(n2397)
         );
  NAND2_X2 U4350 ( .A1(decode_regfile_fpregs_15__17_), .A2(n13263), .ZN(n2398)
         );
  NAND2_X2 U4352 ( .A1(decode_regfile_fpregs_15__16_), .A2(n13262), .ZN(n2399)
         );
  NAND2_X2 U4354 ( .A1(decode_regfile_fpregs_15__15_), .A2(n13262), .ZN(n2400)
         );
  NAND2_X2 U4356 ( .A1(decode_regfile_fpregs_15__14_), .A2(n13263), .ZN(n2401)
         );
  NAND2_X2 U4358 ( .A1(decode_regfile_fpregs_15__13_), .A2(n13262), .ZN(n2402)
         );
  NAND2_X2 U4360 ( .A1(decode_regfile_fpregs_15__12_), .A2(n13262), .ZN(n2403)
         );
  NAND2_X2 U4362 ( .A1(decode_regfile_fpregs_15__11_), .A2(n13263), .ZN(n2404)
         );
  NAND2_X2 U4364 ( .A1(decode_regfile_fpregs_15__10_), .A2(n13262), .ZN(n2405)
         );
  NAND2_X2 U4366 ( .A1(decode_regfile_fpregs_15__0_), .A2(n13263), .ZN(n2406)
         );
  NAND2_X2 U4369 ( .A1(decode_regfile_fpregs_14__9_), .A2(n13257), .ZN(n2409)
         );
  NAND2_X2 U4371 ( .A1(decode_regfile_fpregs_14__8_), .A2(n13259), .ZN(n2410)
         );
  NAND2_X2 U4373 ( .A1(decode_regfile_fpregs_14__7_), .A2(n13259), .ZN(n2411)
         );
  NAND2_X2 U4375 ( .A1(decode_regfile_fpregs_14__6_), .A2(n13259), .ZN(n2412)
         );
  NAND2_X2 U4377 ( .A1(decode_regfile_fpregs_14__5_), .A2(n13259), .ZN(n2413)
         );
  NAND2_X2 U4379 ( .A1(decode_regfile_fpregs_14__4_), .A2(n13259), .ZN(n2414)
         );
  NAND2_X2 U4381 ( .A1(decode_regfile_fpregs_14__3_), .A2(n13259), .ZN(n2415)
         );
  NAND2_X2 U4383 ( .A1(decode_regfile_fpregs_14__31_), .A2(n13259), .ZN(n2416)
         );
  NAND2_X2 U4385 ( .A1(decode_regfile_fpregs_14__30_), .A2(n13258), .ZN(n2417)
         );
  NAND2_X2 U4387 ( .A1(decode_regfile_fpregs_14__2_), .A2(n13258), .ZN(n2418)
         );
  NAND2_X2 U4389 ( .A1(decode_regfile_fpregs_14__29_), .A2(n13258), .ZN(n2419)
         );
  NAND2_X2 U4391 ( .A1(decode_regfile_fpregs_14__28_), .A2(n13258), .ZN(n2420)
         );
  NAND2_X2 U4393 ( .A1(decode_regfile_fpregs_14__27_), .A2(n13258), .ZN(n2421)
         );
  NAND2_X2 U4395 ( .A1(decode_regfile_fpregs_14__26_), .A2(n13258), .ZN(n2422)
         );
  NAND2_X2 U4397 ( .A1(decode_regfile_fpregs_14__25_), .A2(n13258), .ZN(n2423)
         );
  NAND2_X2 U4399 ( .A1(decode_regfile_fpregs_14__24_), .A2(n13258), .ZN(n2424)
         );
  NAND2_X2 U4401 ( .A1(decode_regfile_fpregs_14__23_), .A2(n13258), .ZN(n2425)
         );
  NAND2_X2 U4403 ( .A1(decode_regfile_fpregs_14__22_), .A2(n13258), .ZN(n2426)
         );
  NAND2_X2 U4405 ( .A1(decode_regfile_fpregs_14__21_), .A2(n13258), .ZN(n2427)
         );
  NAND2_X2 U4407 ( .A1(decode_regfile_fpregs_14__20_), .A2(n13258), .ZN(n2428)
         );
  NAND2_X2 U4409 ( .A1(decode_regfile_fpregs_14__1_), .A2(n13258), .ZN(n2429)
         );
  NAND2_X2 U4411 ( .A1(decode_regfile_fpregs_14__19_), .A2(n13258), .ZN(n2430)
         );
  NAND2_X2 U4413 ( .A1(decode_regfile_fpregs_14__18_), .A2(n13258), .ZN(n2431)
         );
  NAND2_X2 U4415 ( .A1(decode_regfile_fpregs_14__17_), .A2(n13258), .ZN(n2432)
         );
  NAND2_X2 U4417 ( .A1(decode_regfile_fpregs_14__16_), .A2(n13257), .ZN(n2433)
         );
  NAND2_X2 U4419 ( .A1(decode_regfile_fpregs_14__15_), .A2(n13257), .ZN(n2434)
         );
  NAND2_X2 U4421 ( .A1(decode_regfile_fpregs_14__14_), .A2(n13258), .ZN(n2435)
         );
  NAND2_X2 U4423 ( .A1(decode_regfile_fpregs_14__13_), .A2(n13257), .ZN(n2436)
         );
  NAND2_X2 U4425 ( .A1(decode_regfile_fpregs_14__12_), .A2(n13257), .ZN(n2437)
         );
  NAND2_X2 U4427 ( .A1(decode_regfile_fpregs_14__11_), .A2(n13258), .ZN(n2438)
         );
  NAND2_X2 U4429 ( .A1(decode_regfile_fpregs_14__10_), .A2(n13257), .ZN(n2439)
         );
  NAND2_X2 U4431 ( .A1(decode_regfile_fpregs_14__0_), .A2(n13258), .ZN(n2440)
         );
  NAND2_X2 U4434 ( .A1(decode_regfile_fpregs_13__9_), .A2(n13252), .ZN(n2442)
         );
  NAND2_X2 U4436 ( .A1(decode_regfile_fpregs_13__8_), .A2(n2441), .ZN(n2443)
         );
  NAND2_X2 U4438 ( .A1(decode_regfile_fpregs_13__7_), .A2(n2441), .ZN(n2444)
         );
  NAND2_X2 U4440 ( .A1(decode_regfile_fpregs_13__6_), .A2(n2441), .ZN(n2445)
         );
  NAND2_X2 U4442 ( .A1(decode_regfile_fpregs_13__5_), .A2(n2441), .ZN(n2446)
         );
  NAND2_X2 U4444 ( .A1(decode_regfile_fpregs_13__4_), .A2(n2441), .ZN(n2447)
         );
  NAND2_X2 U4446 ( .A1(decode_regfile_fpregs_13__3_), .A2(n2441), .ZN(n2448)
         );
  NAND2_X2 U4448 ( .A1(decode_regfile_fpregs_13__31_), .A2(n2441), .ZN(n2449)
         );
  NAND2_X2 U4450 ( .A1(decode_regfile_fpregs_13__30_), .A2(n13253), .ZN(n2450)
         );
  NAND2_X2 U4452 ( .A1(decode_regfile_fpregs_13__2_), .A2(n13253), .ZN(n2451)
         );
  NAND2_X2 U4454 ( .A1(decode_regfile_fpregs_13__29_), .A2(n13253), .ZN(n2452)
         );
  NAND2_X2 U4456 ( .A1(decode_regfile_fpregs_13__28_), .A2(n13253), .ZN(n2453)
         );
  NAND2_X2 U4458 ( .A1(decode_regfile_fpregs_13__27_), .A2(n13253), .ZN(n2454)
         );
  NAND2_X2 U4460 ( .A1(decode_regfile_fpregs_13__26_), .A2(n13253), .ZN(n2455)
         );
  NAND2_X2 U4462 ( .A1(decode_regfile_fpregs_13__25_), .A2(n13253), .ZN(n2456)
         );
  NAND2_X2 U4464 ( .A1(decode_regfile_fpregs_13__24_), .A2(n13253), .ZN(n2457)
         );
  NAND2_X2 U4466 ( .A1(decode_regfile_fpregs_13__23_), .A2(n13253), .ZN(n2458)
         );
  NAND2_X2 U4468 ( .A1(decode_regfile_fpregs_13__22_), .A2(n13253), .ZN(n2459)
         );
  NAND2_X2 U4470 ( .A1(decode_regfile_fpregs_13__21_), .A2(n13253), .ZN(n2460)
         );
  NAND2_X2 U4472 ( .A1(decode_regfile_fpregs_13__20_), .A2(n13253), .ZN(n2461)
         );
  NAND2_X2 U4474 ( .A1(decode_regfile_fpregs_13__1_), .A2(n13253), .ZN(n2462)
         );
  NAND2_X2 U4476 ( .A1(decode_regfile_fpregs_13__19_), .A2(n13253), .ZN(n2463)
         );
  NAND2_X2 U4478 ( .A1(decode_regfile_fpregs_13__18_), .A2(n13253), .ZN(n2464)
         );
  NAND2_X2 U4480 ( .A1(decode_regfile_fpregs_13__17_), .A2(n13253), .ZN(n2465)
         );
  NAND2_X2 U4482 ( .A1(decode_regfile_fpregs_13__16_), .A2(n13252), .ZN(n2466)
         );
  NAND2_X2 U4484 ( .A1(decode_regfile_fpregs_13__15_), .A2(n13252), .ZN(n2467)
         );
  NAND2_X2 U4486 ( .A1(decode_regfile_fpregs_13__14_), .A2(n13253), .ZN(n2468)
         );
  NAND2_X2 U4488 ( .A1(decode_regfile_fpregs_13__13_), .A2(n13252), .ZN(n2469)
         );
  NAND2_X2 U4490 ( .A1(decode_regfile_fpregs_13__12_), .A2(n13252), .ZN(n2470)
         );
  NAND2_X2 U4492 ( .A1(decode_regfile_fpregs_13__11_), .A2(n13253), .ZN(n2471)
         );
  NAND2_X2 U4494 ( .A1(decode_regfile_fpregs_13__10_), .A2(n13252), .ZN(n2472)
         );
  NAND2_X2 U4496 ( .A1(decode_regfile_fpregs_13__0_), .A2(n13253), .ZN(n2473)
         );
  NAND2_X2 U4497 ( .A1(n2407), .A2(n800), .ZN(n2441) );
  NAND2_X2 U4500 ( .A1(decode_regfile_fpregs_12__9_), .A2(n13247), .ZN(n2476)
         );
  NAND2_X2 U4502 ( .A1(decode_regfile_fpregs_12__8_), .A2(n2475), .ZN(n2477)
         );
  NAND2_X2 U4504 ( .A1(decode_regfile_fpregs_12__7_), .A2(n2475), .ZN(n2478)
         );
  NAND2_X2 U4506 ( .A1(decode_regfile_fpregs_12__6_), .A2(n2475), .ZN(n2479)
         );
  NAND2_X2 U4508 ( .A1(decode_regfile_fpregs_12__5_), .A2(n2475), .ZN(n2480)
         );
  NAND2_X2 U4510 ( .A1(decode_regfile_fpregs_12__4_), .A2(n2475), .ZN(n2481)
         );
  NAND2_X2 U4512 ( .A1(decode_regfile_fpregs_12__3_), .A2(n2475), .ZN(n2482)
         );
  NAND2_X2 U4514 ( .A1(decode_regfile_fpregs_12__31_), .A2(n2475), .ZN(n2483)
         );
  NAND2_X2 U4516 ( .A1(decode_regfile_fpregs_12__30_), .A2(n13248), .ZN(n2484)
         );
  NAND2_X2 U4518 ( .A1(decode_regfile_fpregs_12__2_), .A2(n13248), .ZN(n2485)
         );
  NAND2_X2 U4520 ( .A1(decode_regfile_fpregs_12__29_), .A2(n13248), .ZN(n2486)
         );
  NAND2_X2 U4522 ( .A1(decode_regfile_fpregs_12__28_), .A2(n13248), .ZN(n2487)
         );
  NAND2_X2 U4524 ( .A1(decode_regfile_fpregs_12__27_), .A2(n13248), .ZN(n2488)
         );
  NAND2_X2 U4526 ( .A1(decode_regfile_fpregs_12__26_), .A2(n13248), .ZN(n2489)
         );
  NAND2_X2 U4528 ( .A1(decode_regfile_fpregs_12__25_), .A2(n13248), .ZN(n2490)
         );
  NAND2_X2 U4530 ( .A1(decode_regfile_fpregs_12__24_), .A2(n13248), .ZN(n2491)
         );
  NAND2_X2 U4532 ( .A1(decode_regfile_fpregs_12__23_), .A2(n13248), .ZN(n2492)
         );
  NAND2_X2 U4534 ( .A1(decode_regfile_fpregs_12__22_), .A2(n13248), .ZN(n2493)
         );
  NAND2_X2 U4536 ( .A1(decode_regfile_fpregs_12__21_), .A2(n13248), .ZN(n2494)
         );
  NAND2_X2 U4538 ( .A1(decode_regfile_fpregs_12__20_), .A2(n13248), .ZN(n2495)
         );
  NAND2_X2 U4540 ( .A1(decode_regfile_fpregs_12__1_), .A2(n13248), .ZN(n2496)
         );
  NAND2_X2 U4542 ( .A1(decode_regfile_fpregs_12__19_), .A2(n13248), .ZN(n2497)
         );
  NAND2_X2 U4544 ( .A1(decode_regfile_fpregs_12__18_), .A2(n13248), .ZN(n2498)
         );
  NAND2_X2 U4546 ( .A1(decode_regfile_fpregs_12__17_), .A2(n13248), .ZN(n2499)
         );
  NAND2_X2 U4548 ( .A1(decode_regfile_fpregs_12__16_), .A2(n13247), .ZN(n2500)
         );
  NAND2_X2 U4550 ( .A1(decode_regfile_fpregs_12__15_), .A2(n13247), .ZN(n2501)
         );
  NAND2_X2 U4552 ( .A1(decode_regfile_fpregs_12__14_), .A2(n13248), .ZN(n2502)
         );
  NAND2_X2 U4554 ( .A1(decode_regfile_fpregs_12__13_), .A2(n13247), .ZN(n2503)
         );
  NAND2_X2 U4556 ( .A1(decode_regfile_fpregs_12__12_), .A2(n13247), .ZN(n2504)
         );
  NAND2_X2 U4558 ( .A1(decode_regfile_fpregs_12__11_), .A2(n13248), .ZN(n2505)
         );
  NAND2_X2 U4560 ( .A1(decode_regfile_fpregs_12__10_), .A2(n13247), .ZN(n2506)
         );
  NAND2_X2 U4562 ( .A1(decode_regfile_fpregs_12__0_), .A2(n13248), .ZN(n2507)
         );
  NAND2_X2 U4563 ( .A1(n2407), .A2(n834), .ZN(n2475) );
  AND2_X2 U4564 ( .A1(n1738), .A2(n836), .ZN(n2407) );
  NAND2_X2 U4568 ( .A1(decode_regfile_fpregs_11__9_), .A2(n13242), .ZN(n2510)
         );
  NAND2_X2 U4570 ( .A1(decode_regfile_fpregs_11__8_), .A2(n13244), .ZN(n2511)
         );
  NAND2_X2 U4572 ( .A1(decode_regfile_fpregs_11__7_), .A2(n13244), .ZN(n2512)
         );
  NAND2_X2 U4574 ( .A1(decode_regfile_fpregs_11__6_), .A2(n13244), .ZN(n2513)
         );
  NAND2_X2 U4576 ( .A1(decode_regfile_fpregs_11__5_), .A2(n13244), .ZN(n2514)
         );
  NAND2_X2 U4578 ( .A1(decode_regfile_fpregs_11__4_), .A2(n13244), .ZN(n2515)
         );
  NAND2_X2 U4580 ( .A1(decode_regfile_fpregs_11__3_), .A2(n13244), .ZN(n2516)
         );
  NAND2_X2 U4582 ( .A1(decode_regfile_fpregs_11__31_), .A2(n13244), .ZN(n2517)
         );
  NAND2_X2 U4584 ( .A1(decode_regfile_fpregs_11__30_), .A2(n13243), .ZN(n2518)
         );
  NAND2_X2 U4586 ( .A1(decode_regfile_fpregs_11__2_), .A2(n13243), .ZN(n2519)
         );
  NAND2_X2 U4588 ( .A1(decode_regfile_fpregs_11__29_), .A2(n13243), .ZN(n2520)
         );
  NAND2_X2 U4590 ( .A1(decode_regfile_fpregs_11__28_), .A2(n13243), .ZN(n2521)
         );
  NAND2_X2 U4592 ( .A1(decode_regfile_fpregs_11__27_), .A2(n13243), .ZN(n2522)
         );
  NAND2_X2 U4594 ( .A1(decode_regfile_fpregs_11__26_), .A2(n13243), .ZN(n2523)
         );
  NAND2_X2 U4596 ( .A1(decode_regfile_fpregs_11__25_), .A2(n13243), .ZN(n2524)
         );
  NAND2_X2 U4598 ( .A1(decode_regfile_fpregs_11__24_), .A2(n13243), .ZN(n2525)
         );
  NAND2_X2 U4600 ( .A1(decode_regfile_fpregs_11__23_), .A2(n13243), .ZN(n2526)
         );
  NAND2_X2 U4602 ( .A1(decode_regfile_fpregs_11__22_), .A2(n13243), .ZN(n2527)
         );
  NAND2_X2 U4604 ( .A1(decode_regfile_fpregs_11__21_), .A2(n13243), .ZN(n2528)
         );
  NAND2_X2 U4606 ( .A1(decode_regfile_fpregs_11__20_), .A2(n13243), .ZN(n2529)
         );
  NAND2_X2 U4608 ( .A1(decode_regfile_fpregs_11__1_), .A2(n13243), .ZN(n2530)
         );
  NAND2_X2 U4610 ( .A1(decode_regfile_fpregs_11__19_), .A2(n13243), .ZN(n2531)
         );
  NAND2_X2 U4612 ( .A1(decode_regfile_fpregs_11__18_), .A2(n13243), .ZN(n2532)
         );
  NAND2_X2 U4614 ( .A1(decode_regfile_fpregs_11__17_), .A2(n13243), .ZN(n2533)
         );
  NAND2_X2 U4616 ( .A1(decode_regfile_fpregs_11__16_), .A2(n13242), .ZN(n2534)
         );
  NAND2_X2 U4618 ( .A1(decode_regfile_fpregs_11__15_), .A2(n13242), .ZN(n2535)
         );
  NAND2_X2 U4620 ( .A1(decode_regfile_fpregs_11__14_), .A2(n13243), .ZN(n2536)
         );
  NAND2_X2 U4622 ( .A1(decode_regfile_fpregs_11__13_), .A2(n13242), .ZN(n2537)
         );
  NAND2_X2 U4624 ( .A1(decode_regfile_fpregs_11__12_), .A2(n13242), .ZN(n2538)
         );
  NAND2_X2 U4626 ( .A1(decode_regfile_fpregs_11__11_), .A2(n13243), .ZN(n2539)
         );
  NAND2_X2 U4628 ( .A1(decode_regfile_fpregs_11__10_), .A2(n13242), .ZN(n2540)
         );
  NAND2_X2 U4630 ( .A1(decode_regfile_fpregs_11__0_), .A2(n13243), .ZN(n2541)
         );
  NAND2_X2 U4634 ( .A1(decode_regfile_fpregs_10__9_), .A2(n13237), .ZN(n2543)
         );
  NAND2_X2 U4636 ( .A1(decode_regfile_fpregs_10__8_), .A2(n13239), .ZN(n2544)
         );
  NAND2_X2 U4638 ( .A1(decode_regfile_fpregs_10__7_), .A2(n13239), .ZN(n2545)
         );
  NAND2_X2 U4640 ( .A1(decode_regfile_fpregs_10__6_), .A2(n13239), .ZN(n2546)
         );
  NAND2_X2 U4642 ( .A1(decode_regfile_fpregs_10__5_), .A2(n13239), .ZN(n2547)
         );
  NAND2_X2 U4644 ( .A1(decode_regfile_fpregs_10__4_), .A2(n13239), .ZN(n2548)
         );
  NAND2_X2 U4646 ( .A1(decode_regfile_fpregs_10__3_), .A2(n13239), .ZN(n2549)
         );
  NAND2_X2 U4648 ( .A1(decode_regfile_fpregs_10__31_), .A2(n13239), .ZN(n2550)
         );
  NAND2_X2 U4650 ( .A1(decode_regfile_fpregs_10__30_), .A2(n13238), .ZN(n2551)
         );
  NAND2_X2 U4652 ( .A1(decode_regfile_fpregs_10__2_), .A2(n13238), .ZN(n2552)
         );
  NAND2_X2 U4654 ( .A1(decode_regfile_fpregs_10__29_), .A2(n13238), .ZN(n2553)
         );
  NAND2_X2 U4656 ( .A1(decode_regfile_fpregs_10__28_), .A2(n13238), .ZN(n2554)
         );
  NAND2_X2 U4658 ( .A1(decode_regfile_fpregs_10__27_), .A2(n13238), .ZN(n2555)
         );
  NAND2_X2 U4660 ( .A1(decode_regfile_fpregs_10__26_), .A2(n13238), .ZN(n2556)
         );
  NAND2_X2 U4662 ( .A1(decode_regfile_fpregs_10__25_), .A2(n13238), .ZN(n2557)
         );
  NAND2_X2 U4664 ( .A1(decode_regfile_fpregs_10__24_), .A2(n13238), .ZN(n2558)
         );
  NAND2_X2 U4666 ( .A1(decode_regfile_fpregs_10__23_), .A2(n13238), .ZN(n2559)
         );
  NAND2_X2 U4668 ( .A1(decode_regfile_fpregs_10__22_), .A2(n13238), .ZN(n2560)
         );
  NAND2_X2 U4670 ( .A1(decode_regfile_fpregs_10__21_), .A2(n13238), .ZN(n2561)
         );
  NAND2_X2 U4672 ( .A1(decode_regfile_fpregs_10__20_), .A2(n13238), .ZN(n2562)
         );
  NAND2_X2 U4674 ( .A1(decode_regfile_fpregs_10__1_), .A2(n13238), .ZN(n2563)
         );
  NAND2_X2 U4676 ( .A1(decode_regfile_fpregs_10__19_), .A2(n13238), .ZN(n2564)
         );
  NAND2_X2 U4678 ( .A1(decode_regfile_fpregs_10__18_), .A2(n13238), .ZN(n2565)
         );
  NAND2_X2 U4680 ( .A1(decode_regfile_fpregs_10__17_), .A2(n13238), .ZN(n2566)
         );
  NAND2_X2 U4682 ( .A1(decode_regfile_fpregs_10__16_), .A2(n13237), .ZN(n2567)
         );
  NAND2_X2 U4684 ( .A1(decode_regfile_fpregs_10__15_), .A2(n13237), .ZN(n2568)
         );
  NAND2_X2 U4686 ( .A1(decode_regfile_fpregs_10__14_), .A2(n13238), .ZN(n2569)
         );
  NAND2_X2 U4688 ( .A1(decode_regfile_fpregs_10__13_), .A2(n13237), .ZN(n2570)
         );
  NAND2_X2 U4690 ( .A1(decode_regfile_fpregs_10__12_), .A2(n13237), .ZN(n2571)
         );
  NAND2_X2 U4692 ( .A1(decode_regfile_fpregs_10__11_), .A2(n13238), .ZN(n2572)
         );
  NAND2_X2 U4694 ( .A1(decode_regfile_fpregs_10__10_), .A2(n13237), .ZN(n2573)
         );
  NAND2_X2 U4696 ( .A1(decode_regfile_fpregs_10__0_), .A2(n13238), .ZN(n2574)
         );
  AND2_X2 U4700 ( .A1(n1738), .A2(n461), .ZN(n1571) );
  NAND2_X2 U4704 ( .A1(decode_regfile_fpregs_0__9_), .A2(n13232), .ZN(n2576)
         );
  AOI22_X2 U4705 ( .A1(n16357), .A2(decode_regfile_N122), .B1(n16552), .B2(
        n13228), .ZN(n1506) );
  AOI22_X2 U4707 ( .A1(rgwrite_busWout[9]), .A2(n13781), .B1(
        rgwrite_delayslot2out[9]), .B2(n13779), .ZN(n2578) );
  NAND2_X2 U4709 ( .A1(decode_regfile_fpregs_0__8_), .A2(n2575), .ZN(n2580) );
  AOI22_X2 U4710 ( .A1(n16357), .A2(decode_regfile_N123), .B1(n16553), .B2(
        n13229), .ZN(n1509) );
  AOI22_X2 U4712 ( .A1(rgwrite_busWout[8]), .A2(n13781), .B1(
        rgwrite_delayslot2out[8]), .B2(rgwrite_jalout), .ZN(n2581) );
  NAND2_X2 U4714 ( .A1(decode_regfile_fpregs_0__7_), .A2(n2575), .ZN(n2582) );
  AOI22_X2 U4715 ( .A1(n16357), .A2(decode_regfile_N124), .B1(n16554), .B2(
        n13229), .ZN(n1511) );
  AOI22_X2 U4717 ( .A1(rgwrite_busWout[7]), .A2(n13781), .B1(
        rgwrite_delayslot2out[7]), .B2(rgwrite_jalout), .ZN(n2583) );
  NAND2_X2 U4719 ( .A1(decode_regfile_fpregs_0__6_), .A2(n2575), .ZN(n2584) );
  AOI22_X2 U4720 ( .A1(n16357), .A2(decode_regfile_N125), .B1(n16555), .B2(
        n13229), .ZN(n1513) );
  AOI22_X2 U4722 ( .A1(rgwrite_busWout[6]), .A2(n13781), .B1(
        rgwrite_delayslot2out[6]), .B2(rgwrite_jalout), .ZN(n2585) );
  NAND2_X2 U4724 ( .A1(decode_regfile_fpregs_0__5_), .A2(n2575), .ZN(n2586) );
  AOI22_X2 U4725 ( .A1(n16357), .A2(decode_regfile_N126), .B1(n16556), .B2(
        n13229), .ZN(n1515) );
  AOI22_X2 U4727 ( .A1(rgwrite_busWout[5]), .A2(n13781), .B1(
        rgwrite_delayslot2out[5]), .B2(rgwrite_jalout), .ZN(n2587) );
  NAND2_X2 U4729 ( .A1(decode_regfile_fpregs_0__4_), .A2(n2575), .ZN(n2588) );
  AOI22_X2 U4730 ( .A1(n16357), .A2(decode_regfile_N127), .B1(n16557), .B2(
        n13229), .ZN(n1517) );
  AOI22_X2 U4732 ( .A1(rgwrite_busWout[4]), .A2(n13781), .B1(
        rgwrite_delayslot2out[4]), .B2(rgwrite_jalout), .ZN(n2589) );
  NAND2_X2 U4734 ( .A1(decode_regfile_fpregs_0__3_), .A2(n2575), .ZN(n2590) );
  AOI22_X2 U4735 ( .A1(n13128), .A2(decode_regfile_N128), .B1(n16558), .B2(
        n13229), .ZN(n1519) );
  AOI22_X2 U4737 ( .A1(rgwrite_busWout[3]), .A2(n13781), .B1(
        rgwrite_delayslot2out[3]), .B2(rgwrite_jalout), .ZN(n2591) );
  NAND2_X2 U4739 ( .A1(decode_regfile_fpregs_0__31_), .A2(n2575), .ZN(n2592)
         );
  AOI22_X2 U4740 ( .A1(n16357), .A2(decode_regfile_N100), .B1(n16559), .B2(
        n13229), .ZN(n1521) );
  AOI22_X2 U4742 ( .A1(rgwrite_busWout[31]), .A2(n13781), .B1(
        rgwrite_delayslot2out[31]), .B2(rgwrite_jalout), .ZN(n2593) );
  NAND2_X2 U4744 ( .A1(decode_regfile_fpregs_0__30_), .A2(n13233), .ZN(n2594)
         );
  AOI22_X2 U4745 ( .A1(n16357), .A2(decode_regfile_N101), .B1(n16560), .B2(
        n13229), .ZN(n1523) );
  AOI22_X2 U4747 ( .A1(rgwrite_busWout[30]), .A2(n13781), .B1(
        rgwrite_delayslot2out[30]), .B2(rgwrite_jalout), .ZN(n2595) );
  NAND2_X2 U4749 ( .A1(decode_regfile_fpregs_0__2_), .A2(n13233), .ZN(n2596)
         );
  AOI22_X2 U4750 ( .A1(n16357), .A2(decode_regfile_N129), .B1(n16561), .B2(
        n13229), .ZN(n1525) );
  AOI22_X2 U4752 ( .A1(rgwrite_busWout[2]), .A2(n13781), .B1(
        rgwrite_delayslot2out[2]), .B2(rgwrite_jalout), .ZN(n2597) );
  NAND2_X2 U4754 ( .A1(decode_regfile_fpregs_0__29_), .A2(n13233), .ZN(n2598)
         );
  AOI22_X2 U4755 ( .A1(n16357), .A2(decode_regfile_N102), .B1(n16562), .B2(
        n13229), .ZN(n1527) );
  AOI22_X2 U4757 ( .A1(rgwrite_busWout[29]), .A2(n13781), .B1(
        rgwrite_delayslot2out[29]), .B2(n13780), .ZN(n2599) );
  NAND2_X2 U4759 ( .A1(decode_regfile_fpregs_0__28_), .A2(n13233), .ZN(n2600)
         );
  AOI22_X2 U4760 ( .A1(n16357), .A2(decode_regfile_N103), .B1(n16563), .B2(
        n13229), .ZN(n1529) );
  AOI22_X2 U4762 ( .A1(rgwrite_busWout[28]), .A2(n13781), .B1(
        rgwrite_delayslot2out[28]), .B2(n13780), .ZN(n2601) );
  NAND2_X2 U4764 ( .A1(decode_regfile_fpregs_0__27_), .A2(n13233), .ZN(n2602)
         );
  AOI22_X2 U4765 ( .A1(n16357), .A2(decode_regfile_N104), .B1(n16564), .B2(
        n13229), .ZN(n1531) );
  AOI22_X2 U4767 ( .A1(rgwrite_busWout[27]), .A2(n13781), .B1(
        rgwrite_delayslot2out[27]), .B2(n13780), .ZN(n2603) );
  NAND2_X2 U4769 ( .A1(decode_regfile_fpregs_0__26_), .A2(n13233), .ZN(n2604)
         );
  AOI22_X2 U4770 ( .A1(n16357), .A2(decode_regfile_N105), .B1(n16565), .B2(
        n13229), .ZN(n1533) );
  AOI22_X2 U4772 ( .A1(rgwrite_busWout[26]), .A2(n13781), .B1(
        rgwrite_delayslot2out[26]), .B2(n13780), .ZN(n2605) );
  NAND2_X2 U4774 ( .A1(decode_regfile_fpregs_0__25_), .A2(n13233), .ZN(n2606)
         );
  AOI22_X2 U4775 ( .A1(n16357), .A2(decode_regfile_N106), .B1(n16566), .B2(
        n13229), .ZN(n1535) );
  AOI22_X2 U4777 ( .A1(rgwrite_busWout[25]), .A2(n13781), .B1(
        rgwrite_delayslot2out[25]), .B2(n13780), .ZN(n2607) );
  NAND2_X2 U4779 ( .A1(decode_regfile_fpregs_0__24_), .A2(n13233), .ZN(n2608)
         );
  AOI22_X2 U4780 ( .A1(n16357), .A2(decode_regfile_N107), .B1(n16567), .B2(
        n13229), .ZN(n1537) );
  AOI22_X2 U4782 ( .A1(rgwrite_busWout[24]), .A2(n13781), .B1(
        rgwrite_delayslot2out[24]), .B2(n13780), .ZN(n2609) );
  NAND2_X2 U4784 ( .A1(decode_regfile_fpregs_0__23_), .A2(n13233), .ZN(n2610)
         );
  AOI22_X2 U4785 ( .A1(n13128), .A2(decode_regfile_N108), .B1(n16568), .B2(
        n13229), .ZN(n1539) );
  AOI22_X2 U4787 ( .A1(rgwrite_busWout[23]), .A2(n13781), .B1(
        rgwrite_delayslot2out[23]), .B2(n13780), .ZN(n2611) );
  NAND2_X2 U4789 ( .A1(decode_regfile_fpregs_0__22_), .A2(n13233), .ZN(n2612)
         );
  AOI22_X2 U4790 ( .A1(n13128), .A2(decode_regfile_N109), .B1(n16569), .B2(
        n13228), .ZN(n1541) );
  AOI22_X2 U4792 ( .A1(rgwrite_busWout[22]), .A2(n13781), .B1(
        rgwrite_delayslot2out[22]), .B2(n13780), .ZN(n2613) );
  NAND2_X2 U4794 ( .A1(decode_regfile_fpregs_0__21_), .A2(n13233), .ZN(n2614)
         );
  AOI22_X2 U4795 ( .A1(n13128), .A2(decode_regfile_N110), .B1(n16570), .B2(
        n13228), .ZN(n1543) );
  AOI22_X2 U4797 ( .A1(rgwrite_busWout[21]), .A2(n13781), .B1(
        rgwrite_delayslot2out[21]), .B2(n13780), .ZN(n2615) );
  NAND2_X2 U4799 ( .A1(decode_regfile_fpregs_0__20_), .A2(n13233), .ZN(n2616)
         );
  AOI22_X2 U4800 ( .A1(n13128), .A2(decode_regfile_N111), .B1(n16571), .B2(
        n13228), .ZN(n1545) );
  AOI22_X2 U4802 ( .A1(rgwrite_busWout[20]), .A2(n13781), .B1(
        rgwrite_delayslot2out[20]), .B2(n13780), .ZN(n2617) );
  NAND2_X2 U4804 ( .A1(decode_regfile_fpregs_0__1_), .A2(n13233), .ZN(n2618)
         );
  AOI22_X2 U4805 ( .A1(n13128), .A2(decode_regfile_N130), .B1(n16572), .B2(
        n13228), .ZN(n1547) );
  AOI22_X2 U4807 ( .A1(rgwrite_busWout[1]), .A2(n8721), .B1(
        rgwrite_delayslot2out[1]), .B2(n13780), .ZN(n2619) );
  NAND2_X2 U4809 ( .A1(decode_regfile_fpregs_0__19_), .A2(n13233), .ZN(n2620)
         );
  AOI22_X2 U4810 ( .A1(n13128), .A2(decode_regfile_N112), .B1(n16255), .B2(
        n13228), .ZN(n1549) );
  AOI22_X2 U4812 ( .A1(rgwrite_busWout[19]), .A2(n8721), .B1(
        rgwrite_delayslot2out[19]), .B2(n13779), .ZN(n2621) );
  NAND2_X2 U4814 ( .A1(decode_regfile_fpregs_0__18_), .A2(n13233), .ZN(n2622)
         );
  AOI22_X2 U4815 ( .A1(n13128), .A2(decode_regfile_N113), .B1(n16573), .B2(
        n13228), .ZN(n1551) );
  AOI22_X2 U4817 ( .A1(rgwrite_busWout[18]), .A2(n8721), .B1(
        rgwrite_delayslot2out[18]), .B2(n13779), .ZN(n2623) );
  NAND2_X2 U4819 ( .A1(decode_regfile_fpregs_0__17_), .A2(n13233), .ZN(n2624)
         );
  AOI22_X2 U4820 ( .A1(n13128), .A2(decode_regfile_N114), .B1(n16574), .B2(
        n13228), .ZN(n1553) );
  AOI22_X2 U4822 ( .A1(rgwrite_busWout[17]), .A2(n8721), .B1(
        rgwrite_delayslot2out[17]), .B2(n13779), .ZN(n2625) );
  NAND2_X2 U4824 ( .A1(decode_regfile_fpregs_0__16_), .A2(n13232), .ZN(n2626)
         );
  AOI22_X2 U4825 ( .A1(n13128), .A2(decode_regfile_N115), .B1(n16575), .B2(
        n13228), .ZN(n1555) );
  AOI22_X2 U4827 ( .A1(rgwrite_busWout[16]), .A2(n8721), .B1(n13779), .B2(
        rgwrite_delayslot2out[16]), .ZN(n2627) );
  NAND2_X2 U4829 ( .A1(decode_regfile_fpregs_0__15_), .A2(n13232), .ZN(n2628)
         );
  AOI22_X2 U4830 ( .A1(n13128), .A2(decode_regfile_N116), .B1(n16576), .B2(
        n13228), .ZN(n1557) );
  AOI22_X2 U4832 ( .A1(rgwrite_busWout[15]), .A2(n8721), .B1(
        rgwrite_delayslot2out[15]), .B2(n13779), .ZN(n2629) );
  NAND2_X2 U4834 ( .A1(decode_regfile_fpregs_0__14_), .A2(n13233), .ZN(n2630)
         );
  AOI22_X2 U4835 ( .A1(n13128), .A2(decode_regfile_N117), .B1(n16577), .B2(
        n13228), .ZN(n1559) );
  AOI22_X2 U4837 ( .A1(rgwrite_busWout[14]), .A2(n8721), .B1(
        rgwrite_delayslot2out[14]), .B2(n13779), .ZN(n2631) );
  NAND2_X2 U4839 ( .A1(decode_regfile_fpregs_0__13_), .A2(n13232), .ZN(n2632)
         );
  AOI22_X2 U4840 ( .A1(n13128), .A2(decode_regfile_N118), .B1(n16578), .B2(
        n13228), .ZN(n1561) );
  AOI22_X2 U4842 ( .A1(rgwrite_busWout[13]), .A2(n8721), .B1(
        rgwrite_delayslot2out[13]), .B2(n13779), .ZN(n2633) );
  NAND2_X2 U4844 ( .A1(decode_regfile_fpregs_0__12_), .A2(n13232), .ZN(n2634)
         );
  AOI22_X2 U4845 ( .A1(n13128), .A2(decode_regfile_N119), .B1(n16579), .B2(
        n13228), .ZN(n1563) );
  AOI22_X2 U4847 ( .A1(rgwrite_busWout[12]), .A2(n8721), .B1(
        rgwrite_delayslot2out[12]), .B2(n13779), .ZN(n2635) );
  NAND2_X2 U4849 ( .A1(decode_regfile_fpregs_0__11_), .A2(n13233), .ZN(n2636)
         );
  AOI22_X2 U4850 ( .A1(n13128), .A2(decode_regfile_N120), .B1(n16580), .B2(
        n13228), .ZN(n1565) );
  AOI22_X2 U4852 ( .A1(rgwrite_busWout[11]), .A2(n8721), .B1(
        rgwrite_delayslot2out[11]), .B2(n13779), .ZN(n2637) );
  NAND2_X2 U4854 ( .A1(decode_regfile_fpregs_0__10_), .A2(n13232), .ZN(n2638)
         );
  AOI22_X2 U4855 ( .A1(n13128), .A2(decode_regfile_N121), .B1(n16581), .B2(
        n13228), .ZN(n1567) );
  AOI22_X2 U4857 ( .A1(rgwrite_busWout[10]), .A2(n8721), .B1(
        rgwrite_delayslot2out[10]), .B2(n13779), .ZN(n2639) );
  NAND2_X2 U4859 ( .A1(decode_regfile_fpregs_0__0_), .A2(n13233), .ZN(n2640)
         );
  NAND2_X2 U4860 ( .A1(n1772), .A2(n834), .ZN(n2575) );
  AND2_X2 U4862 ( .A1(n1738), .A2(n664), .ZN(n1772) );
  AOI22_X2 U4866 ( .A1(n16357), .A2(decode_regfile_N131), .B1(n16582), .B2(
        n13228), .ZN(n1569) );
  AOI22_X2 U4869 ( .A1(rgwrite_busWout[0]), .A2(n8721), .B1(
        rgwrite_delayslot2out[0]), .B2(n13780), .ZN(n2641) );
  NAND2_X2 U4872 ( .A1(fpoint_3[0]), .A2(n8724), .ZN(n267) );
  NAND4_X2 U4874 ( .A1(n281), .A2(n280), .A3(n302), .A4(n2642), .ZN(
        decode_decoder_N279) );
  OAI221_X2 U4877 ( .B1(imm32_0[1]), .B2(n2645), .C1(n2646), .C2(n2647), .A(
        n2648), .ZN(n2643) );
  NAND4_X2 U4878 ( .A1(n2649), .A2(n292), .A3(n301), .A4(n2650), .ZN(
        decode_decoder_N278) );
  OAI22_X2 U4883 ( .A1(n2655), .A2(n2646), .B1(n2647), .B2(imm32_0[1]), .ZN(
        n2654) );
  NAND2_X2 U4884 ( .A1(n2656), .A2(n148), .ZN(n2648) );
  NAND2_X2 U4885 ( .A1(n2646), .A2(n202), .ZN(n148) );
  AOI22_X2 U4891 ( .A1(n8726), .A2(n16586), .B1(n2665), .B2(n2657), .ZN(n2663)
         );
  NAND4_X2 U4893 ( .A1(n2666), .A2(n281), .A3(n302), .A4(n2667), .ZN(
        decode_decoder_N276) );
  NAND4_X2 U4896 ( .A1(n16584), .A2(n2672), .A3(n2673), .A4(n2652), .ZN(n2668)
         );
  NAND2_X2 U4902 ( .A1(imm32_0[2]), .A2(n8750), .ZN(n147) );
  NAND2_X2 U4903 ( .A1(n2658), .A2(n16586), .ZN(n2672) );
  OAI22_X2 U4908 ( .A1(imm32_0[1]), .A2(n2655), .B1(n202), .B2(n2645), .ZN(
        n2662) );
  NAND2_X2 U4910 ( .A1(n8726), .A2(n8748), .ZN(n202) );
  NAND2_X2 U4915 ( .A1(imm32_0[5]), .A2(n8749), .ZN(n2675) );
  NAND4_X2 U4920 ( .A1(n8728), .A2(n8751), .A3(n2677), .A4(n8707), .ZN(n137)
         );
  NAND2_X2 U4925 ( .A1(n305), .A2(n16598), .ZN(decode_decoder_N275) );
  NOR4_X2 U4927 ( .A1(n284), .A2(n309), .A3(n16593), .A4(n2678), .ZN(n305) );
  NAND4_X2 U4928 ( .A1(n280), .A2(n281), .A3(n282), .A4(n293), .ZN(n2678) );
  NAND4_X2 U4929 ( .A1(instruction_1[28]), .A2(n2679), .A3(n16596), .A4(n8741), 
        .ZN(n293) );
  NAND2_X2 U4930 ( .A1(n2681), .A2(n16599), .ZN(n282) );
  NAND2_X2 U4931 ( .A1(n16603), .A2(n2683), .ZN(n281) );
  NAND2_X2 U4936 ( .A1(n296), .A2(n16603), .ZN(n301) );
  OAI211_X2 U4937 ( .C1(n2690), .C2(n2691), .A(n2692), .B(n143), .ZN(n2669) );
  NAND2_X2 U4940 ( .A1(n16603), .A2(n2685), .ZN(n292) );
  OAI211_X2 U4946 ( .C1(n2683), .C2(n16596), .A(n2697), .B(instruction_1[31]), 
        .ZN(n2692) );
  OAI211_X2 U4949 ( .C1(n2689), .C2(n2695), .A(n2666), .B(n2649), .ZN(n306) );
  NAND2_X2 U4954 ( .A1(n16604), .A2(n296), .ZN(n277) );
  NAND2_X2 U4955 ( .A1(n16604), .A2(n2685), .ZN(n283) );
  NAND2_X2 U4969 ( .A1(n2699), .A2(n163), .ZN(decode_decoder_N274) );
  AND2_X2 U4971 ( .A1(n2686), .A2(n8742), .ZN(n2681) );
  NAND2_X2 U4977 ( .A1(n2699), .A2(n149), .ZN(n160) );
  AND2_X2 U4978 ( .A1(n220), .A2(n2700), .ZN(n2699) );
  NAND2_X2 U4981 ( .A1(instruction_1[27]), .A2(n8716), .ZN(n2689) );
  NAND4_X2 U4989 ( .A1(n2701), .A2(n2702), .A3(n2703), .A4(n2704), .ZN(
        aluout_0[9]) );
  XOR2_X2 U4997 ( .A(n16331), .B(n2729), .Z(n2723) );
  NAND4_X2 U4999 ( .A1(n2735), .A2(n2736), .A3(n2737), .A4(n2738), .ZN(
        aluout_0[8]) );
  AOI221_X2 U5000 ( .B1(n2739), .B2(n2740), .C1(n16347), .C2(n2742), .A(n2743), 
        .ZN(n2738) );
  OAI22_X2 U5001 ( .A1(n2744), .A2(n13220), .B1(n2745), .B2(n2746), .ZN(n2743)
         );
  XOR2_X2 U5007 ( .A(n2755), .B(n2756), .Z(n2754) );
  NAND4_X2 U5009 ( .A1(n2762), .A2(n2763), .A3(n2764), .A4(n2765), .ZN(
        aluout_0[7]) );
  AOI221_X2 U5010 ( .B1(n2766), .B2(n2767), .C1(n16350), .C2(n2769), .A(n2770), 
        .ZN(n2765) );
  OAI22_X2 U5011 ( .A1(n2771), .A2(n2772), .B1(n2773), .B2(n13220), .ZN(n2770)
         );
  AOI221_X2 U5015 ( .B1(n13114), .B2(n2779), .C1(n2733), .C2(n2780), .A(n2781), 
        .ZN(n2763) );
  OAI22_X2 U5016 ( .A1(n13784), .A2(n2783), .B1(n2784), .B2(n2785), .ZN(n2781)
         );
  XNOR2_X2 U5017 ( .A(n2786), .B(n2787), .ZN(n2783) );
  NAND4_X2 U5019 ( .A1(n2792), .A2(n2793), .A3(n2794), .A4(n2795), .ZN(
        aluout_0[6]) );
  AOI221_X2 U5020 ( .B1(n2796), .B2(n2797), .C1(n16353), .C2(n2799), .A(n2800), 
        .ZN(n2795) );
  OAI22_X2 U5021 ( .A1(n2801), .A2(n2772), .B1(n2802), .B2(n13220), .ZN(n2800)
         );
  AOI221_X2 U5026 ( .B1(n13114), .B2(n2808), .C1(n2733), .C2(n2809), .A(n2810), 
        .ZN(n2793) );
  OAI22_X2 U5027 ( .A1(n13784), .A2(n2811), .B1(n16513), .B2(n2785), .ZN(n2810) );
  XOR2_X2 U5028 ( .A(n2813), .B(n2814), .Z(n2811) );
  NAND4_X2 U5030 ( .A1(n2818), .A2(n2819), .A3(n2820), .A4(n2821), .ZN(
        aluout_0[5]) );
  AOI221_X2 U5031 ( .B1(n2822), .B2(n2823), .C1(n16447), .C2(n2825), .A(n2826), 
        .ZN(n2821) );
  OAI22_X2 U5032 ( .A1(n2827), .A2(n2772), .B1(n2828), .B2(n13220), .ZN(n2826)
         );
  AOI221_X2 U5036 ( .B1(n13114), .B2(n2831), .C1(n2733), .C2(n2832), .A(n2833), 
        .ZN(n2819) );
  OAI22_X2 U5037 ( .A1(n13784), .A2(n2834), .B1(n16488), .B2(n2785), .ZN(n2833) );
  XNOR2_X2 U5038 ( .A(n2836), .B(n2837), .ZN(n2834) );
  NAND4_X2 U5041 ( .A1(n2841), .A2(n2842), .A3(n2843), .A4(n2844), .ZN(
        aluout_0[4]) );
  OAI22_X2 U5047 ( .A1(n13227), .A2(n2845), .B1(n16551), .B2(n2856), .ZN(n2853) );
  XOR2_X2 U5049 ( .A(n2858), .B(n2859), .Z(n2857) );
  AOI22_X2 U5050 ( .A1(n16458), .A2(n16469), .B1(n16548), .B2(n16451), .ZN(
        n2841) );
  NAND4_X2 U5052 ( .A1(n16463), .A2(n2863), .A3(n2864), .A4(n2865), .ZN(
        aluout_0[3]) );
  AOI221_X2 U5055 ( .B1(n8696), .B2(n2777), .C1(n16469), .C2(n2778), .A(n2872), 
        .ZN(n2870) );
  OAI22_X2 U5056 ( .A1(n2771), .A2(n2873), .B1(n2874), .B2(n13103), .ZN(n2872)
         );
  AOI221_X2 U5057 ( .B1(n13183), .B2(n13119), .C1(n13171), .C2(n8651), .A(
        n2878), .ZN(n2874) );
  OAI22_X2 U5058 ( .A1(n13197), .A2(n2880), .B1(n13196), .B2(n2882), .ZN(n2878) );
  AOI221_X2 U5059 ( .B1(n8648), .B2(n13183), .C1(n13115), .C2(n13171), .A(
        n2883), .ZN(n2771) );
  OAI22_X2 U5060 ( .A1(n2884), .A2(n13196), .B1(n2885), .B2(n13197), .ZN(n2883) );
  AOI22_X2 U5062 ( .A1(n13218), .A2(n2887), .B1(n2888), .B2(execstage_ALU_N160), .ZN(n2864) );
  XOR2_X2 U5063 ( .A(n16479), .B(n2890), .Z(n2888) );
  OAI22_X2 U5066 ( .A1(n2895), .A2(n2721), .B1(n2896), .B2(n2897), .ZN(n2894)
         );
  OAI211_X2 U5067 ( .C1(n2898), .C2(n8744), .A(n2900), .B(n2901), .ZN(
        aluout_0[31]) );
  OAI221_X2 U5073 ( .B1(n2917), .B2(n13194), .C1(n8737), .C2(n13184), .A(n2920), .ZN(n2907) );
  XOR2_X2 U5075 ( .A(n2923), .B(n2924), .Z(n2903) );
  XOR2_X2 U5076 ( .A(n2925), .B(n2902), .Z(n2924) );
  XOR2_X2 U5078 ( .A(n13132), .B(n2929), .Z(n2923) );
  NAND2_X2 U5079 ( .A1(execstage_BusA[30]), .A2(n2930), .ZN(n2929) );
  AOI22_X2 U5080 ( .A1(n2931), .A2(n2932), .B1(n16438), .B2(n2934), .ZN(n2900)
         );
  XNOR2_X2 U5083 ( .A(n2935), .B(n2936), .ZN(n2931) );
  XOR2_X2 U5084 ( .A(n2937), .B(n2938), .Z(n2936) );
  XOR2_X2 U5085 ( .A(n2939), .B(n2940), .Z(n2938) );
  XOR2_X2 U5086 ( .A(n2941), .B(n2942), .Z(n2940) );
  XOR2_X2 U5087 ( .A(n2943), .B(n2944), .Z(n2942) );
  XNOR2_X2 U5090 ( .A(n2950), .B(n2951), .ZN(n2941) );
  OAI22_X2 U5092 ( .A1(n2955), .A2(n2956), .B1(n2957), .B2(n2958), .ZN(n2950)
         );
  XOR2_X2 U5093 ( .A(n2959), .B(n2960), .Z(n2939) );
  XOR2_X2 U5094 ( .A(n2961), .B(n2962), .Z(n2960) );
  AND2_X2 U5096 ( .A1(n2965), .A2(n2966), .ZN(n2961) );
  XOR2_X2 U5097 ( .A(n2967), .B(n2968), .Z(n2959) );
  XOR2_X2 U5099 ( .A(n2971), .B(n2972), .Z(n2967) );
  XOR2_X2 U5100 ( .A(n2973), .B(n2974), .Z(n2972) );
  XOR2_X2 U5101 ( .A(n2975), .B(n2976), .Z(n2974) );
  XOR2_X2 U5105 ( .A(n2982), .B(n2983), .Z(n2973) );
  NAND2_X2 U5106 ( .A1(n16433), .A2(n13115), .ZN(n2983) );
  XOR2_X2 U5108 ( .A(n2988), .B(n2989), .Z(n2971) );
  XOR2_X2 U5109 ( .A(n2990), .B(n2991), .Z(n2989) );
  XOR2_X2 U5110 ( .A(n2992), .B(n2993), .Z(n2991) );
  XOR2_X2 U5111 ( .A(n2994), .B(n2995), .Z(n2993) );
  XNOR2_X2 U5112 ( .A(n2996), .B(n2997), .ZN(n2995) );
  XOR2_X2 U5116 ( .A(n3005), .B(n3006), .Z(n2992) );
  XOR2_X2 U5117 ( .A(n3007), .B(n3008), .Z(n3006) );
  XOR2_X2 U5118 ( .A(n3009), .B(n3010), .Z(n3008) );
  XOR2_X2 U5119 ( .A(n3011), .B(n3012), .Z(n3010) );
  XOR2_X2 U5120 ( .A(n3013), .B(n3014), .Z(n3012) );
  XOR2_X2 U5121 ( .A(n3015), .B(n3016), .Z(n3014) );
  XOR2_X2 U5122 ( .A(n3017), .B(n3018), .Z(n3016) );
  XOR2_X2 U5123 ( .A(n3019), .B(n3020), .Z(n3018) );
  XOR2_X2 U5124 ( .A(n3021), .B(n3022), .Z(n3020) );
  XOR2_X2 U5125 ( .A(n3023), .B(n3024), .Z(n3022) );
  XOR2_X2 U5126 ( .A(n3025), .B(n3026), .Z(n3024) );
  AND2_X2 U5127 ( .A1(n3027), .A2(n3028), .ZN(n3026) );
  NAND2_X2 U5128 ( .A1(n3029), .A2(n16257), .ZN(n3025) );
  XOR2_X2 U5129 ( .A(n3031), .B(n3032), .Z(n3023) );
  XOR2_X2 U5130 ( .A(n3033), .B(n3034), .Z(n3032) );
  NAND2_X2 U5131 ( .A1(n13113), .A2(execstage_BusA[14]), .ZN(n3034) );
  NAND2_X2 U5133 ( .A1(execstage_BusA[19]), .A2(n13164), .ZN(n3031) );
  XOR2_X2 U5134 ( .A(n3040), .B(n3041), .Z(n3021) );
  XOR2_X2 U5135 ( .A(n3042), .B(n3043), .Z(n3041) );
  XOR2_X2 U5136 ( .A(n3044), .B(n3045), .Z(n3043) );
  XOR2_X2 U5137 ( .A(n3046), .B(n3047), .Z(n3045) );
  NAND2_X2 U5139 ( .A1(n3050), .A2(n16334), .ZN(n3046) );
  XOR2_X2 U5140 ( .A(n3052), .B(n3053), .Z(n3044) );
  XOR2_X2 U5141 ( .A(n3054), .B(n3055), .Z(n3053) );
  XOR2_X2 U5142 ( .A(n3056), .B(n3057), .Z(n3055) );
  NAND2_X2 U5143 ( .A1(execstage_BusA[27]), .A2(n13192), .ZN(n3057) );
  NAND2_X2 U5144 ( .A1(execstage_BusA[22]), .A2(n13158), .ZN(n3056) );
  XOR2_X2 U5145 ( .A(n3058), .B(n3059), .Z(n3054) );
  XOR2_X2 U5148 ( .A(n3066), .B(n3067), .Z(n3052) );
  XOR2_X2 U5149 ( .A(n3068), .B(n3069), .Z(n3067) );
  AND2_X2 U5151 ( .A1(n3072), .A2(n3073), .ZN(n3068) );
  XOR2_X2 U5152 ( .A(n3074), .B(n3075), .Z(n3066) );
  XOR2_X2 U5154 ( .A(n3077), .B(n3078), .Z(n3074) );
  XOR2_X2 U5155 ( .A(n3079), .B(n3080), .Z(n3078) );
  XOR2_X2 U5156 ( .A(n3081), .B(n3082), .Z(n3080) );
  NAND2_X2 U5158 ( .A1(n3085), .A2(n2921), .ZN(n3081) );
  XOR2_X2 U5159 ( .A(n3086), .B(n3087), .Z(n3079) );
  AOI22_X2 U5160 ( .A1(n3088), .A2(n3089), .B1(n3090), .B2(n3091), .ZN(n3087)
         );
  NAND2_X2 U5161 ( .A1(execstage_BusA[29]), .A2(n13177), .ZN(n3086) );
  XOR2_X2 U5162 ( .A(n3093), .B(n3094), .Z(n3077) );
  XOR2_X2 U5163 ( .A(n3095), .B(n3096), .Z(n3094) );
  NAND2_X2 U5164 ( .A1(execstage_BusA[28]), .A2(n13204), .ZN(n3096) );
  NAND2_X2 U5165 ( .A1(execstage_BusA[26]), .A2(n13207), .ZN(n3095) );
  XOR2_X2 U5166 ( .A(n3097), .B(n3098), .Z(n3093) );
  OAI221_X2 U5168 ( .B1(execstage_ALU_ra_row2_31_), .B2(n3101), .C1(n13186), 
        .C2(n8658), .A(n3103), .ZN(n3097) );
  NAND2_X2 U5170 ( .A1(execstage_BusA[30]), .A2(n13199), .ZN(n3101) );
  XOR2_X2 U5171 ( .A(n3105), .B(n3106), .Z(n3042) );
  XOR2_X2 U5172 ( .A(n3107), .B(n3108), .Z(n3106) );
  NAND2_X2 U5173 ( .A1(n3109), .A2(n3110), .ZN(n3108) );
  NAND2_X2 U5174 ( .A1(execstage_BusA[23]), .A2(n13217), .ZN(n3107) );
  XOR2_X2 U5175 ( .A(n3111), .B(n3112), .Z(n3105) );
  NAND2_X2 U5176 ( .A1(execstage_BusA[18]), .A2(n13166), .ZN(n3112) );
  NAND2_X2 U5178 ( .A1(n3117), .A2(n3118), .ZN(n3040) );
  XOR2_X2 U5179 ( .A(n3119), .B(n3120), .Z(n3019) );
  XNOR2_X2 U5180 ( .A(n3121), .B(n3122), .ZN(n3120) );
  XOR2_X2 U5183 ( .A(n3128), .B(n3129), .Z(n3119) );
  NAND2_X2 U5185 ( .A1(execstage_BusA[25]), .A2(n13211), .ZN(n3128) );
  NAND2_X2 U5186 ( .A1(n3132), .A2(n3133), .ZN(n3017) );
  XOR2_X2 U5187 ( .A(n3134), .B(n3135), .Z(n3015) );
  XOR2_X2 U5188 ( .A(n3136), .B(n3137), .Z(n3135) );
  XOR2_X2 U5189 ( .A(n3138), .B(n3139), .Z(n3137) );
  NAND2_X2 U5190 ( .A1(n16406), .A2(n13122), .ZN(n3139) );
  XOR2_X2 U5193 ( .A(n3146), .B(n3147), .Z(n3134) );
  NAND2_X2 U5195 ( .A1(n3150), .A2(n3151), .ZN(n3146) );
  XOR2_X2 U5196 ( .A(n3152), .B(n3153), .Z(n3013) );
  XOR2_X2 U5197 ( .A(n3154), .B(n3155), .Z(n3153) );
  NAND2_X2 U5198 ( .A1(execstage_BusA[21]), .A2(n13161), .ZN(n3155) );
  NAND2_X2 U5199 ( .A1(execstage_BusA[16]), .A2(n13168), .ZN(n3154) );
  XNOR2_X2 U5200 ( .A(n3158), .B(n3159), .ZN(n3152) );
  NAND2_X2 U5203 ( .A1(n3165), .A2(n3166), .ZN(n3011) );
  XOR2_X2 U5204 ( .A(n3167), .B(n3168), .Z(n3009) );
  XOR2_X2 U5205 ( .A(n3169), .B(n3170), .Z(n3168) );
  XOR2_X2 U5206 ( .A(n3171), .B(n3172), .Z(n3170) );
  NAND2_X2 U5207 ( .A1(n16435), .A2(n13116), .ZN(n3172) );
  XOR2_X2 U5210 ( .A(n3179), .B(n3180), .Z(n3167) );
  NAND2_X2 U5212 ( .A1(n3183), .A2(n3184), .ZN(n3179) );
  XOR2_X2 U5213 ( .A(n3185), .B(n3186), .Z(n3007) );
  XOR2_X2 U5214 ( .A(n3187), .B(n3188), .Z(n3186) );
  NAND2_X2 U5215 ( .A1(execstage_BusA[17]), .A2(n13179), .ZN(n3188) );
  NAND2_X2 U5216 ( .A1(n13112), .A2(execstage_BusA[12]), .ZN(n3187) );
  XNOR2_X2 U5217 ( .A(n3191), .B(n3192), .ZN(n3185) );
  XOR2_X2 U5220 ( .A(n3198), .B(n3199), .Z(n3005) );
  NAND2_X2 U5222 ( .A1(n3202), .A2(n3203), .ZN(n3198) );
  NAND2_X2 U5223 ( .A1(n3204), .A2(n3205), .ZN(n2990) );
  XOR2_X2 U5224 ( .A(n3206), .B(n3207), .Z(n2988) );
  NAND2_X2 U5226 ( .A1(n13111), .A2(n13118), .ZN(n3206) );
  XOR2_X2 U5228 ( .A(n3213), .B(n3214), .Z(n2935) );
  XOR2_X2 U5229 ( .A(n3215), .B(n3216), .Z(n3214) );
  NAND2_X2 U5230 ( .A1(n16426), .A2(n13791), .ZN(n3216) );
  NAND2_X2 U5231 ( .A1(n16437), .A2(execstage_BusA[1]), .ZN(n3215) );
  NAND2_X2 U5232 ( .A1(n3218), .A2(n3219), .ZN(n3213) );
  AOI221_X2 U5233 ( .B1(n3220), .B2(n13171), .C1(n16438), .C2(n16548), .A(
        n3221), .ZN(n2898) );
  NAND2_X2 U5234 ( .A1(n3222), .A2(n13219), .ZN(n3221) );
  AOI221_X2 U5236 ( .B1(n16549), .B2(n3226), .C1(n13130), .C2(n3227), .A(n3228), .ZN(n3225) );
  OAI222_X2 U5238 ( .A1(n3230), .A2(n3231), .B1(n13192), .B2(n3232), .C1(
        n16467), .C2(n13190), .ZN(n3226) );
  NAND2_X2 U5243 ( .A1(n3242), .A2(n3243), .ZN(n3239) );
  AOI22_X2 U5246 ( .A1(n16437), .A2(n3248), .B1(n3249), .B2(execstage_ALU_N160), .ZN(n3223) );
  XOR2_X2 U5247 ( .A(n2927), .B(n2926), .Z(n3249) );
  AOI22_X2 U5248 ( .A1(n3250), .A2(execstage_BusA[29]), .B1(n3251), .B2(n3252), 
        .ZN(n2926) );
  XOR2_X2 U5249 ( .A(n8658), .B(n2930), .Z(n2927) );
  XOR2_X2 U5250 ( .A(execstage_ALU_sel), .B(n16437), .Z(n2930) );
  OAI221_X2 U5251 ( .B1(n3212), .B2(n13226), .C1(n2896), .C2(n8658), .A(n13219), .ZN(n3248) );
  XOR2_X2 U5252 ( .A(n2956), .B(n2955), .Z(n3212) );
  XNOR2_X2 U5253 ( .A(n2958), .B(n2957), .ZN(n2955) );
  XNOR2_X2 U5254 ( .A(n3219), .B(n3218), .ZN(n2957) );
  XOR2_X2 U5255 ( .A(n2963), .B(n2964), .Z(n3218) );
  NAND2_X2 U5256 ( .A1(n16426), .A2(execstage_BusA[2]), .ZN(n2964) );
  NAND2_X2 U5258 ( .A1(n3253), .A2(n3254), .ZN(n2949) );
  XOR2_X2 U5260 ( .A(n2948), .B(n2947), .Z(n3253) );
  XNOR2_X2 U5261 ( .A(n2965), .B(n2966), .ZN(n2947) );
  XOR2_X2 U5262 ( .A(n2977), .B(n2978), .Z(n2966) );
  NAND2_X2 U5263 ( .A1(n16429), .A2(execstage_BusA[4]), .ZN(n2978) );
  NAND2_X2 U5265 ( .A1(n3259), .A2(n3260), .ZN(n2954) );
  XOR2_X2 U5267 ( .A(n2952), .B(n2953), .Z(n3259) );
  XOR2_X2 U5268 ( .A(n2981), .B(n2980), .Z(n2953) );
  XNOR2_X2 U5269 ( .A(n2998), .B(n2999), .ZN(n2980) );
  NAND2_X2 U5270 ( .A1(n16433), .A2(execstage_BusA[6]), .ZN(n2999) );
  NAND2_X2 U5272 ( .A1(n3264), .A2(n3265), .ZN(n2987) );
  XOR2_X2 U5274 ( .A(n2986), .B(n2985), .Z(n3264) );
  XNOR2_X2 U5275 ( .A(n3205), .B(n3204), .ZN(n2985) );
  XOR2_X2 U5276 ( .A(n3181), .B(n3182), .Z(n3204) );
  NAND2_X2 U5277 ( .A1(n13111), .A2(execstage_BusA[8]), .ZN(n3182) );
  NAND2_X2 U5279 ( .A1(n3269), .A2(n3270), .ZN(n3176) );
  XOR2_X2 U5281 ( .A(n3175), .B(n3174), .Z(n3269) );
  XNOR2_X2 U5282 ( .A(n3184), .B(n3183), .ZN(n3174) );
  XOR2_X2 U5283 ( .A(n3193), .B(n3194), .Z(n3183) );
  NAND2_X2 U5284 ( .A1(n16409), .A2(n8694), .ZN(n3194) );
  NAND2_X2 U5286 ( .A1(n3275), .A2(n3276), .ZN(n3002) );
  XOR2_X2 U5288 ( .A(n3000), .B(n3001), .Z(n3275) );
  XNOR2_X2 U5289 ( .A(n3203), .B(n3202), .ZN(n3001) );
  XOR2_X2 U5290 ( .A(n3148), .B(n3149), .Z(n3202) );
  NAND2_X2 U5291 ( .A1(n13109), .A2(execstage_BusA[12]), .ZN(n3149) );
  NAND2_X2 U5293 ( .A1(n3281), .A2(n3282), .ZN(n3143) );
  XOR2_X2 U5295 ( .A(n3142), .B(n3141), .Z(n3281) );
  XNOR2_X2 U5296 ( .A(n3151), .B(n3150), .ZN(n3141) );
  XOR2_X2 U5297 ( .A(n3160), .B(n3161), .Z(n3150) );
  NAND2_X2 U5298 ( .A1(n13107), .A2(execstage_BusA[14]), .ZN(n3161) );
  NAND2_X2 U5300 ( .A1(n3287), .A2(n3288), .ZN(n3197) );
  XOR2_X2 U5302 ( .A(n3196), .B(n3195), .Z(n3287) );
  XNOR2_X2 U5303 ( .A(n3166), .B(n3165), .ZN(n3195) );
  XOR2_X2 U5304 ( .A(n16257), .B(n3029), .Z(n3165) );
  NAND2_X2 U5308 ( .A1(n3295), .A2(n3296), .ZN(n3038) );
  XOR2_X2 U5311 ( .A(n3037), .B(n3036), .Z(n3295) );
  XNOR2_X2 U5312 ( .A(n3027), .B(n3028), .ZN(n3036) );
  XOR2_X2 U5313 ( .A(n3123), .B(n3124), .Z(n3028) );
  NAND2_X2 U5314 ( .A1(execstage_BusA[18]), .A2(n13164), .ZN(n3124) );
  NAND2_X2 U5316 ( .A1(n3301), .A2(n3302), .ZN(n3164) );
  XOR2_X2 U5318 ( .A(n3162), .B(n3163), .Z(n3301) );
  XNOR2_X2 U5319 ( .A(n3133), .B(n3132), .ZN(n3163) );
  XOR2_X2 U5320 ( .A(n3048), .B(n3049), .Z(n3132) );
  NAND2_X2 U5321 ( .A1(execstage_BusA[20]), .A2(n13161), .ZN(n3049) );
  NAND2_X2 U5323 ( .A1(n3306), .A2(n3307), .ZN(n3116) );
  XOR2_X2 U5326 ( .A(n3115), .B(n3114), .Z(n3306) );
  XNOR2_X2 U5327 ( .A(n3110), .B(n3109), .ZN(n3114) );
  XOR2_X2 U5328 ( .A(n16334), .B(n3050), .Z(n3109) );
  NAND2_X2 U5332 ( .A1(n3314), .A2(n3315), .ZN(n3127) );
  XOR2_X2 U5335 ( .A(n3125), .B(n3126), .Z(n3314) );
  XNOR2_X2 U5336 ( .A(n3118), .B(n3117), .ZN(n3126) );
  XOR2_X2 U5337 ( .A(n3070), .B(n3071), .Z(n3117) );
  NAND2_X2 U5338 ( .A1(execstage_BusA[24]), .A2(n13211), .ZN(n3071) );
  NAND2_X2 U5340 ( .A1(n3320), .A2(n3321), .ZN(n3065) );
  XOR2_X2 U5343 ( .A(n3064), .B(n3063), .Z(n3320) );
  XNOR2_X2 U5344 ( .A(n3072), .B(n3073), .ZN(n3063) );
  XNOR2_X2 U5345 ( .A(n3083), .B(n3326), .ZN(n3073) );
  NAND2_X2 U5348 ( .A1(n3327), .A2(n3328), .ZN(n3062) );
  XOR2_X2 U5350 ( .A(n3061), .B(n3060), .Z(n3327) );
  XNOR2_X2 U5351 ( .A(n3089), .B(n3088), .ZN(n3060) );
  XOR2_X2 U5352 ( .A(n3090), .B(n3091), .Z(n3088) );
  XOR2_X2 U5353 ( .A(n3100), .B(n3099), .Z(n3091) );
  XNOR2_X2 U5357 ( .A(n3085), .B(n2921), .ZN(n3100) );
  NAND2_X2 U5361 ( .A1(execstage_BusA[27]), .A2(n13204), .ZN(n3061) );
  NAND2_X2 U5364 ( .A1(execstage_BusA[25]), .A2(n13207), .ZN(n3064) );
  NAND2_X2 U5367 ( .A1(execstage_BusA[23]), .A2(n13214), .ZN(n3125) );
  NAND2_X2 U5370 ( .A1(execstage_BusA[21]), .A2(n13158), .ZN(n3115) );
  NAND2_X2 U5373 ( .A1(execstage_BusA[19]), .A2(n13182), .ZN(n3162) );
  NAND2_X2 U5375 ( .A1(execstage_BusA[17]), .A2(n13166), .ZN(n3037) );
  NAND2_X2 U5379 ( .A1(n13113), .A2(n8655), .ZN(n3142) );
  NAND2_X2 U5381 ( .A1(n13112), .A2(n8652), .ZN(n3000) );
  NAND2_X2 U5383 ( .A1(n16406), .A2(n8648), .ZN(n3175) );
  NAND2_X2 U5385 ( .A1(n16431), .A2(n13115), .ZN(n2986) );
  NAND2_X2 U5387 ( .A1(n16435), .A2(n13119), .ZN(n2952) );
  NAND2_X2 U5389 ( .A1(n16427), .A2(n13791), .ZN(n2948) );
  NAND2_X2 U5391 ( .A1(n16424), .A2(execstage_BusA[1]), .ZN(n2958) );
  AOI221_X2 U5394 ( .B1(n3394), .B2(n13783), .C1(n13114), .C2(n3395), .A(n3396), .ZN(n3393) );
  OAI221_X2 U5395 ( .B1(n3397), .B2(n3398), .C1(n3399), .C2(n13174), .A(n3400), 
        .ZN(n3396) );
  OAI211_X2 U5396 ( .C1(n3401), .C2(n16464), .A(n3403), .B(n13190), .ZN(n3400)
         );
  AOI22_X2 U5398 ( .A1(n2807), .A2(n16469), .B1(n2806), .B2(n8696), .ZN(n3404)
         );
  OAI22_X2 U5399 ( .A1(n2801), .A2(n2873), .B1(n3405), .B2(n13103), .ZN(n3401)
         );
  AOI221_X2 U5400 ( .B1(n16545), .B2(n13194), .C1(n13183), .C2(
        execstage_BusA[4]), .A(n3407), .ZN(n3405) );
  AOI221_X2 U5402 ( .B1(execstage_BusA[8]), .B2(n13187), .C1(n13116), .C2(
        n13171), .A(n3410), .ZN(n2801) );
  OAI22_X2 U5403 ( .A1(n3411), .A2(n13196), .B1(n3412), .B2(n13198), .ZN(n3410) );
  XOR2_X2 U5406 ( .A(n3416), .B(n3417), .Z(n3394) );
  AOI22_X2 U5408 ( .A1(n16548), .A2(n3421), .B1(n13218), .B2(execstage_BusA[2]), .ZN(n3391) );
  OAI22_X2 U5411 ( .A1(n16420), .A2(n2721), .B1(n3428), .B2(n3429), .ZN(n3425)
         );
  OAI221_X2 U5413 ( .B1(n13186), .B2(n8713), .C1(n13169), .C2(n8737), .A(n3435), .ZN(n3432) );
  AOI22_X2 U5414 ( .A1(n16528), .A2(n13198), .B1(n16524), .B2(n13195), .ZN(
        n3435) );
  AOI22_X2 U5421 ( .A1(n16424), .A2(n3446), .B1(n3447), .B2(execstage_ALU_N160), .ZN(n3422) );
  XOR2_X2 U5422 ( .A(n3251), .B(n3252), .Z(n3447) );
  XOR2_X2 U5423 ( .A(execstage_BusA[29]), .B(n3250), .Z(n3252) );
  XNOR2_X2 U5424 ( .A(n13132), .B(n16424), .ZN(n3250) );
  OAI22_X2 U5425 ( .A1(n16425), .A2(n8735), .B1(n3449), .B2(n3450), .ZN(n3251)
         );
  OAI221_X2 U5427 ( .B1(n13227), .B2(n3390), .C1(n2896), .C2(n8737), .A(n13220), .ZN(n3446) );
  XOR2_X2 U5428 ( .A(n3386), .B(n3387), .Z(n3390) );
  NAND2_X2 U5430 ( .A1(n3388), .A2(n3453), .ZN(n3386) );
  OR3_X2 U5432 ( .A1(n3455), .A2(n13152), .A3(n3456), .ZN(n3388) );
  NAND2_X2 U5434 ( .A1(n3457), .A2(n3458), .ZN(n3257) );
  XOR2_X2 U5436 ( .A(n3256), .B(n3255), .Z(n3457) );
  XNOR2_X2 U5437 ( .A(n3383), .B(n3382), .ZN(n3255) );
  NAND2_X2 U5439 ( .A1(n3384), .A2(n3465), .ZN(n3383) );
  OR3_X2 U5441 ( .A1(n2946), .A2(n13790), .A3(n3467), .ZN(n3384) );
  XNOR2_X2 U5442 ( .A(n3262), .B(n16181), .ZN(n3467) );
  NAND2_X2 U5446 ( .A1(n3263), .A2(n3473), .ZN(n3262) );
  OR3_X2 U5448 ( .A1(n3474), .A2(n8738), .A3(n3475), .ZN(n3263) );
  XNOR2_X2 U5449 ( .A(n3380), .B(n3379), .ZN(n3475) );
  NAND2_X2 U5451 ( .A1(n3381), .A2(n3479), .ZN(n3380) );
  OR3_X2 U5453 ( .A1(n3480), .A2(n13143), .A3(n3481), .ZN(n3381) );
  XNOR2_X2 U5454 ( .A(n3267), .B(n16184), .ZN(n3481) );
  NAND2_X2 U5457 ( .A1(n3268), .A2(n3486), .ZN(n3267) );
  OR3_X2 U5459 ( .A1(n3004), .A2(n8715), .A3(n3488), .ZN(n3268) );
  XNOR2_X2 U5460 ( .A(n3376), .B(n3375), .ZN(n3488) );
  NAND2_X2 U5462 ( .A1(n3377), .A2(n3492), .ZN(n3376) );
  OR3_X2 U5464 ( .A1(n3494), .A2(n8739), .A3(n3495), .ZN(n3377) );
  XNOR2_X2 U5465 ( .A(n3272), .B(n3271), .ZN(n3495) );
  NAND2_X2 U5467 ( .A1(n3273), .A2(n3499), .ZN(n3272) );
  OR3_X2 U5469 ( .A1(n3500), .A2(n8714), .A3(n3501), .ZN(n3273) );
  XNOR2_X2 U5470 ( .A(n3373), .B(n16185), .ZN(n3501) );
  NAND2_X2 U5473 ( .A1(n3374), .A2(n3506), .ZN(n3373) );
  OR3_X2 U5475 ( .A1(n3178), .A2(n13146), .A3(n3508), .ZN(n3374) );
  XNOR2_X2 U5476 ( .A(n3278), .B(n16186), .ZN(n3508) );
  NAND2_X2 U5479 ( .A1(n3279), .A2(n3513), .ZN(n3278) );
  OR3_X2 U5481 ( .A1(n3515), .A2(n13136), .A3(n3516), .ZN(n3279) );
  XNOR2_X2 U5482 ( .A(n3370), .B(n16187), .ZN(n3516) );
  NAND2_X2 U5485 ( .A1(n3371), .A2(n3521), .ZN(n3370) );
  OR3_X2 U5487 ( .A1(n13110), .A2(n8736), .A3(n3522), .ZN(n3371) );
  XNOR2_X2 U5488 ( .A(n3284), .B(n16188), .ZN(n3522) );
  NAND2_X2 U5491 ( .A1(n3285), .A2(n3527), .ZN(n3284) );
  OR3_X2 U5493 ( .A1(n3529), .A2(n8695), .A3(n3530), .ZN(n3285) );
  XNOR2_X2 U5494 ( .A(n3367), .B(n16258), .ZN(n3530) );
  NAND2_X2 U5497 ( .A1(n3368), .A2(n3535), .ZN(n3367) );
  OR3_X2 U5499 ( .A1(n3145), .A2(n8710), .A3(n3536), .ZN(n3368) );
  XNOR2_X2 U5500 ( .A(n3290), .B(n16259), .ZN(n3536) );
  NAND2_X2 U5503 ( .A1(n3291), .A2(n3541), .ZN(n3290) );
  OR3_X2 U5505 ( .A1(n3543), .A2(n8657), .A3(n3544), .ZN(n3291) );
  XOR2_X2 U5506 ( .A(n3365), .B(n3363), .Z(n3544) );
  NAND2_X2 U5507 ( .A1(n3364), .A2(n3545), .ZN(n3363) );
  OR3_X2 U5509 ( .A1(n8645), .A2(n13178), .A3(n3546), .ZN(n3364) );
  XOR2_X2 U5510 ( .A(n3300), .B(n3298), .Z(n3546) );
  NAND2_X2 U5511 ( .A1(n3299), .A2(n3547), .ZN(n3298) );
  OR3_X2 U5513 ( .A1(n8734), .A2(n13165), .A3(n3549), .ZN(n3299) );
  XNOR2_X2 U5514 ( .A(n3360), .B(n16262), .ZN(n3549) );
  NAND2_X2 U5517 ( .A1(n3361), .A2(n3554), .ZN(n3360) );
  OR3_X2 U5519 ( .A1(n8647), .A2(n13162), .A3(n3557), .ZN(n3361) );
  XNOR2_X2 U5520 ( .A(n3304), .B(n3303), .ZN(n3557) );
  NAND2_X2 U5522 ( .A1(n3305), .A2(n3561), .ZN(n3304) );
  OR3_X2 U5524 ( .A1(n8650), .A2(n3130), .A3(n3563), .ZN(n3305) );
  XOR2_X2 U5525 ( .A(n3357), .B(n3355), .Z(n3563) );
  NAND2_X2 U5526 ( .A1(n3356), .A2(n3564), .ZN(n3355) );
  OR3_X2 U5528 ( .A1(n8654), .A2(n13159), .A3(n3567), .ZN(n3356) );
  XOR2_X2 U5529 ( .A(n3311), .B(n3309), .Z(n3567) );
  NAND2_X2 U5530 ( .A1(n3310), .A2(n3568), .ZN(n3309) );
  OR3_X2 U5532 ( .A1(n8730), .A2(n13157), .A3(n3570), .ZN(n3310) );
  XOR2_X2 U5533 ( .A(n3353), .B(n3351), .Z(n3570) );
  NAND2_X2 U5534 ( .A1(n3352), .A2(n3571), .ZN(n3351) );
  OR3_X2 U5536 ( .A1(n8646), .A2(n13215), .A3(n3573), .ZN(n3352) );
  XOR2_X2 U5537 ( .A(n3319), .B(n3317), .Z(n3573) );
  NAND2_X2 U5538 ( .A1(n3318), .A2(n3574), .ZN(n3317) );
  OR3_X2 U5540 ( .A1(n8653), .A2(n13212), .A3(n3575), .ZN(n3318) );
  XOR2_X2 U5541 ( .A(n3349), .B(n3347), .Z(n3575) );
  NAND2_X2 U5542 ( .A1(n3348), .A2(n3576), .ZN(n3347) );
  OR3_X2 U5544 ( .A1(n8656), .A2(n13209), .A3(n3578), .ZN(n3348) );
  XOR2_X2 U5545 ( .A(n3325), .B(n3323), .Z(n3578) );
  NAND2_X2 U5546 ( .A1(n3324), .A2(n3579), .ZN(n3323) );
  OR3_X2 U5548 ( .A1(n8731), .A2(n13205), .A3(n3580), .ZN(n3324) );
  XOR2_X2 U5549 ( .A(n3345), .B(n3343), .Z(n3580) );
  XOR2_X2 U5552 ( .A(n16375), .B(n3330), .Z(n3582) );
  NAND2_X2 U5553 ( .A1(n3331), .A2(n3583), .ZN(n3330) );
  OR3_X2 U5555 ( .A1(n8733), .A2(n13201), .A3(n3584), .ZN(n3331) );
  XNOR2_X2 U5556 ( .A(n3340), .B(n16379), .ZN(n3584) );
  NAND2_X2 U5560 ( .A1(n3341), .A2(n3590), .ZN(n3340) );
  OR3_X2 U5562 ( .A1(n8713), .A2(n13175), .A3(n3591), .ZN(n3341) );
  XOR2_X2 U5563 ( .A(n3332), .B(n3336), .Z(n3591) );
  NAND2_X2 U5581 ( .A1(n16427), .A2(n13792), .ZN(n3256) );
  AOI221_X2 U5583 ( .B1(n16549), .B2(n3631), .C1(n13131), .C2(n3632), .A(n3633), .ZN(n3630) );
  OAI222_X2 U5586 ( .A1(n13192), .A2(n3634), .B1(n3635), .B2(n13189), .C1(
        n3636), .C2(n3231), .ZN(n3631) );
  OAI22_X2 U5589 ( .A1(n13170), .A2(n8735), .B1(n13198), .B2(n3641), .ZN(n3637) );
  AOI22_X2 U5597 ( .A1(n16426), .A2(n3654), .B1(n3655), .B2(execstage_ALU_N160), .ZN(n3628) );
  XOR2_X2 U5598 ( .A(n3450), .B(n3449), .Z(n3655) );
  AOI22_X2 U5599 ( .A1(n3656), .A2(execstage_BusA[27]), .B1(n3657), .B2(n3658), 
        .ZN(n3449) );
  XOR2_X2 U5600 ( .A(n8735), .B(n3451), .Z(n3450) );
  XNOR2_X2 U5601 ( .A(n13132), .B(n16426), .ZN(n3451) );
  OAI221_X2 U5602 ( .B1(n13227), .B2(n3452), .C1(n2896), .C2(n8735), .A(n13220), .ZN(n3654) );
  XOR2_X2 U5603 ( .A(n3460), .B(n3459), .Z(n3452) );
  NAND2_X2 U5605 ( .A1(n3461), .A2(n3660), .ZN(n3460) );
  OR3_X2 U5607 ( .A1(n3209), .A2(n13152), .A3(n3661), .ZN(n3461) );
  XNOR2_X2 U5608 ( .A(n3463), .B(n3462), .ZN(n3661) );
  AND3_X2 U5612 ( .A1(n16429), .A2(n13792), .A3(n3666), .ZN(n3464) );
  XNOR2_X2 U5613 ( .A(n3472), .B(n3470), .ZN(n3666) );
  NAND2_X2 U5614 ( .A1(n3471), .A2(n3667), .ZN(n3470) );
  OR3_X2 U5616 ( .A1(n3474), .A2(n13790), .A3(n3668), .ZN(n3471) );
  XNOR2_X2 U5617 ( .A(n3477), .B(n3476), .ZN(n3668) );
  AND3_X2 U5621 ( .A1(n16433), .A2(execstage_BusA[4]), .A3(n3673), .ZN(n3478)
         );
  XOR2_X2 U5622 ( .A(n3484), .B(n3483), .Z(n3673) );
  NAND2_X2 U5624 ( .A1(n3485), .A2(n3677), .ZN(n3484) );
  OR3_X2 U5626 ( .A1(n3004), .A2(n13143), .A3(n3678), .ZN(n3485) );
  XNOR2_X2 U5627 ( .A(n3490), .B(n3489), .ZN(n3678) );
  AND3_X2 U5631 ( .A1(n13111), .A2(n13116), .A3(n3683), .ZN(n3491) );
  XOR2_X2 U5632 ( .A(n3497), .B(n3496), .Z(n3683) );
  AND3_X2 U5636 ( .A1(n16406), .A2(n13115), .A3(n3688), .ZN(n3498) );
  XOR2_X2 U5637 ( .A(n3504), .B(n3503), .Z(n3688) );
  NAND2_X2 U5639 ( .A1(n3505), .A2(n3692), .ZN(n3504) );
  OR3_X2 U5641 ( .A1(n3178), .A2(n8714), .A3(n3693), .ZN(n3505) );
  XNOR2_X2 U5642 ( .A(n3511), .B(n3510), .ZN(n3693) );
  NAND2_X2 U5644 ( .A1(n3512), .A2(n3697), .ZN(n3511) );
  OR3_X2 U5646 ( .A1(n3515), .A2(n13146), .A3(n3698), .ZN(n3512) );
  XNOR2_X2 U5647 ( .A(n3519), .B(n3518), .ZN(n3698) );
  NAND2_X2 U5649 ( .A1(n3520), .A2(n3702), .ZN(n3519) );
  OR3_X2 U5651 ( .A1(n13110), .A2(n13136), .A3(n3703), .ZN(n3520) );
  XNOR2_X2 U5652 ( .A(n3525), .B(n3524), .ZN(n3703) );
  NAND2_X2 U5654 ( .A1(n3526), .A2(n3707), .ZN(n3525) );
  OR3_X2 U5656 ( .A1(n3529), .A2(n8736), .A3(n3708), .ZN(n3526) );
  XNOR2_X2 U5657 ( .A(n3533), .B(n3532), .ZN(n3708) );
  NAND2_X2 U5659 ( .A1(n3534), .A2(n3712), .ZN(n3533) );
  OR3_X2 U5661 ( .A1(n3145), .A2(n8695), .A3(n3713), .ZN(n3534) );
  XNOR2_X2 U5662 ( .A(n3539), .B(n3538), .ZN(n3713) );
  NAND2_X2 U5664 ( .A1(n3540), .A2(n3717), .ZN(n3539) );
  OR3_X2 U5666 ( .A1(n3543), .A2(n8710), .A3(n3718), .ZN(n3540) );
  NAND2_X2 U5668 ( .A1(n3719), .A2(n3720), .ZN(n3627) );
  XOR2_X2 U5670 ( .A(n3625), .B(n3626), .Z(n3719) );
  XNOR2_X2 U5671 ( .A(n3623), .B(n3622), .ZN(n3626) );
  NAND2_X2 U5673 ( .A1(n3624), .A2(n3727), .ZN(n3623) );
  OR3_X2 U5675 ( .A1(n8645), .A2(n13165), .A3(n3728), .ZN(n3624) );
  XNOR2_X2 U5676 ( .A(n3552), .B(n3551), .ZN(n3728) );
  NAND2_X2 U5678 ( .A1(n3553), .A2(n3732), .ZN(n3552) );
  OR3_X2 U5680 ( .A1(n8734), .A2(n13162), .A3(n3733), .ZN(n3553) );
  XNOR2_X2 U5681 ( .A(n3559), .B(n3558), .ZN(n3733) );
  AND3_X2 U5685 ( .A1(execstage_BusA[17]), .A2(n13182), .A3(n3738), .ZN(n3560)
         );
  XOR2_X2 U5686 ( .A(n3619), .B(n3620), .Z(n3738) );
  NAND2_X2 U5687 ( .A1(n3621), .A2(n3739), .ZN(n3620) );
  OR3_X2 U5689 ( .A1(n8650), .A2(n13159), .A3(n3740), .ZN(n3621) );
  XNOR2_X2 U5690 ( .A(n3616), .B(n3617), .ZN(n3740) );
  NAND2_X2 U5691 ( .A1(n3618), .A2(n3741), .ZN(n3617) );
  OR3_X2 U5693 ( .A1(n8654), .A2(n13157), .A3(n3742), .ZN(n3618) );
  XNOR2_X2 U5694 ( .A(n3613), .B(n3614), .ZN(n3742) );
  NAND2_X2 U5695 ( .A1(n3615), .A2(n3743), .ZN(n3614) );
  OR3_X2 U5697 ( .A1(n8730), .A2(n13215), .A3(n3744), .ZN(n3615) );
  XNOR2_X2 U5698 ( .A(n3610), .B(n3611), .ZN(n3744) );
  NAND2_X2 U5699 ( .A1(n3612), .A2(n3745), .ZN(n3611) );
  OR3_X2 U5701 ( .A1(n8646), .A2(n13212), .A3(n3746), .ZN(n3612) );
  XNOR2_X2 U5702 ( .A(n3607), .B(n3608), .ZN(n3746) );
  NAND2_X2 U5703 ( .A1(n3609), .A2(n3747), .ZN(n3608) );
  OR3_X2 U5705 ( .A1(n8653), .A2(n13209), .A3(n3748), .ZN(n3609) );
  XNOR2_X2 U5706 ( .A(n3604), .B(n3605), .ZN(n3748) );
  NAND2_X2 U5707 ( .A1(n3606), .A2(n3749), .ZN(n3605) );
  OR3_X2 U5709 ( .A1(n8656), .A2(n13205), .A3(n3750), .ZN(n3606) );
  XNOR2_X2 U5710 ( .A(n3601), .B(n3602), .ZN(n3750) );
  NAND2_X2 U5711 ( .A1(n3603), .A2(n3751), .ZN(n3602) );
  OR3_X2 U5713 ( .A1(n8731), .A2(n13190), .A3(n3752), .ZN(n3603) );
  XOR2_X2 U5714 ( .A(n3599), .B(n3597), .Z(n3752) );
  NAND2_X2 U5715 ( .A1(n3598), .A2(n3753), .ZN(n3597) );
  OR3_X2 U5717 ( .A1(n8732), .A2(n13201), .A3(n3754), .ZN(n3598) );
  XOR2_X2 U5718 ( .A(n3589), .B(n3587), .Z(n3754) );
  NAND2_X2 U5719 ( .A1(n3588), .A2(n3755), .ZN(n3587) );
  OR3_X2 U5721 ( .A1(n8733), .A2(n13175), .A3(n3756), .ZN(n3588) );
  NAND2_X2 U5723 ( .A1(n3757), .A2(n3758), .ZN(n3594) );
  XOR2_X2 U5726 ( .A(n3593), .B(n2917), .Z(n3757) );
  NAND2_X2 U5727 ( .A1(execstage_BusA[27]), .A2(n13199), .ZN(n3593) );
  NAND4_X2 U5738 ( .A1(n3793), .A2(n3794), .A3(n3795), .A4(n3796), .ZN(
        aluout_0[27]) );
  AOI22_X2 U5742 ( .A1(n3803), .A2(n3244), .B1(n3804), .B2(n16453), .ZN(n3802)
         );
  AND2_X2 U5743 ( .A1(n3806), .A2(n8659), .ZN(n3244) );
  OAI221_X2 U5746 ( .B1(n13227), .B2(n3659), .C1(n2896), .C2(n8713), .A(n13220), .ZN(n3810) );
  XOR2_X2 U5747 ( .A(n3663), .B(n3662), .Z(n3659) );
  NAND2_X2 U5749 ( .A1(n3664), .A2(n3812), .ZN(n3663) );
  OR3_X2 U5751 ( .A1(n2946), .A2(n13152), .A3(n3813), .ZN(n3664) );
  NAND2_X2 U5753 ( .A1(n3814), .A2(n3815), .ZN(n3792) );
  XOR2_X2 U5755 ( .A(n3791), .B(n3790), .Z(n3814) );
  XNOR2_X2 U5756 ( .A(n3670), .B(n3669), .ZN(n3790) );
  NAND2_X2 U5758 ( .A1(n3671), .A2(n3822), .ZN(n3670) );
  OR3_X2 U5760 ( .A1(n3480), .A2(n13790), .A3(n3823), .ZN(n3671) );
  XNOR2_X2 U5761 ( .A(n3675), .B(n3674), .ZN(n3823) );
  AND3_X2 U5766 ( .A1(n16431), .A2(execstage_BusA[4]), .A3(n3829), .ZN(n3676)
         );
  XOR2_X2 U5767 ( .A(n3680), .B(n3679), .Z(n3829) );
  NAND2_X2 U5769 ( .A1(n3681), .A2(n3833), .ZN(n3680) );
  OR3_X2 U5771 ( .A1(n3494), .A2(n13143), .A3(n3834), .ZN(n3681) );
  XNOR2_X2 U5772 ( .A(n3685), .B(n3684), .ZN(n3834) );
  NAND2_X2 U5774 ( .A1(n3686), .A2(n3838), .ZN(n3685) );
  OR3_X2 U5776 ( .A1(n3500), .A2(n8715), .A3(n3839), .ZN(n3686) );
  XNOR2_X2 U5777 ( .A(n3690), .B(n3689), .ZN(n3839) );
  AND3_X2 U5781 ( .A1(n16409), .A2(n13115), .A3(n3844), .ZN(n3691) );
  XOR2_X2 U5782 ( .A(n3695), .B(n3694), .Z(n3844) );
  AND3_X2 U5786 ( .A1(n13112), .A2(execstage_BusA[8]), .A3(n3849), .ZN(n3696)
         );
  XOR2_X2 U5787 ( .A(n3700), .B(n3699), .Z(n3849) );
  AND3_X2 U5791 ( .A1(n13109), .A2(n13118), .A3(n3854), .ZN(n3701) );
  XOR2_X2 U5792 ( .A(n3705), .B(n3704), .Z(n3854) );
  AND3_X2 U5796 ( .A1(n13113), .A2(n13122), .A3(n3859), .ZN(n3706) );
  XOR2_X2 U5797 ( .A(n3710), .B(n3709), .Z(n3859) );
  AND3_X2 U5801 ( .A1(n13107), .A2(n13121), .A3(n3864), .ZN(n3711) );
  XOR2_X2 U5802 ( .A(n3715), .B(n3714), .Z(n3864) );
  AND3_X2 U5806 ( .A1(n13168), .A2(execstage_BusA[12]), .A3(n3869), .ZN(n3716)
         );
  XOR2_X2 U5807 ( .A(n3722), .B(n16265), .Z(n3869) );
  NAND2_X2 U5810 ( .A1(n3723), .A2(n3874), .ZN(n3722) );
  OR3_X2 U5812 ( .A1(n13178), .A2(n8710), .A3(n3875), .ZN(n3723) );
  XNOR2_X2 U5813 ( .A(n3724), .B(n3725), .ZN(n3875) );
  AND3_X2 U5816 ( .A1(execstage_BusA[14]), .A2(n13166), .A3(n3877), .ZN(n3726)
         );
  XOR2_X2 U5817 ( .A(n3730), .B(n3729), .Z(n3877) );
  AND3_X2 U5821 ( .A1(execstage_BusA[15]), .A2(n13164), .A3(n3882), .ZN(n3731)
         );
  XOR2_X2 U5822 ( .A(n3735), .B(n3734), .Z(n3882) );
  NAND2_X2 U5824 ( .A1(n3736), .A2(n3886), .ZN(n3735) );
  OR3_X2 U5826 ( .A1(n8734), .A2(n3130), .A3(n3887), .ZN(n3736) );
  XNOR2_X2 U5827 ( .A(n3787), .B(n3788), .ZN(n3887) );
  AND3_X2 U5830 ( .A1(execstage_BusA[17]), .A2(n13161), .A3(n3889), .ZN(n3789)
         );
  XOR2_X2 U5831 ( .A(n3784), .B(n3785), .Z(n3889) );
  AND3_X2 U5834 ( .A1(execstage_BusA[18]), .A2(n13158), .A3(n3891), .ZN(n3786)
         );
  XOR2_X2 U5835 ( .A(n3781), .B(n3782), .Z(n3891) );
  AND3_X2 U5838 ( .A1(execstage_BusA[19]), .A2(n13217), .A3(n3893), .ZN(n3783)
         );
  XOR2_X2 U5839 ( .A(n3778), .B(n3779), .Z(n3893) );
  AND3_X2 U5842 ( .A1(execstage_BusA[20]), .A2(n13214), .A3(n3895), .ZN(n3780)
         );
  XOR2_X2 U5843 ( .A(n3775), .B(n3776), .Z(n3895) );
  AND3_X2 U5846 ( .A1(execstage_BusA[21]), .A2(n13211), .A3(n3897), .ZN(n3777)
         );
  XOR2_X2 U5847 ( .A(n3772), .B(n3773), .Z(n3897) );
  AND3_X2 U5850 ( .A1(execstage_BusA[22]), .A2(n13208), .A3(n3899), .ZN(n3774)
         );
  XOR2_X2 U5851 ( .A(n3769), .B(n3770), .Z(n3899) );
  AND3_X2 U5854 ( .A1(execstage_BusA[23]), .A2(n13188), .A3(n3901), .ZN(n3771)
         );
  XOR2_X2 U5855 ( .A(n3766), .B(n3767), .Z(n3901) );
  NAND2_X2 U5856 ( .A1(n3768), .A2(n3902), .ZN(n3767) );
  OR3_X2 U5858 ( .A1(n8731), .A2(n13201), .A3(n3903), .ZN(n3768) );
  XNOR2_X2 U5859 ( .A(n3763), .B(n3764), .ZN(n3903) );
  NAND2_X2 U5860 ( .A1(n3765), .A2(n3904), .ZN(n3764) );
  OR3_X2 U5862 ( .A1(n8732), .A2(n13175), .A3(n3905), .ZN(n3765) );
  XOR2_X2 U5863 ( .A(n3762), .B(n3760), .Z(n3905) );
  NAND2_X2 U5864 ( .A1(n3761), .A2(n3906), .ZN(n3760) );
  NAND2_X2 U5866 ( .A1(n16508), .A2(execstage_BusA[26]), .ZN(n3761) );
  NAND2_X2 U5879 ( .A1(n16435), .A2(n13792), .ZN(n3791) );
  OAI222_X2 U5880 ( .A1(n2784), .A2(n13104), .B1(n16496), .B2(n13103), .C1(
        n16495), .C2(n2873), .ZN(n3809) );
  OAI221_X2 U5882 ( .B1(n13186), .B2(n8732), .C1(n13170), .C2(n8713), .A(n3947), .ZN(n2915) );
  AOI22_X2 U5883 ( .A1(n16528), .A2(n13196), .B1(n16527), .B2(n13200), .ZN(
        n3947) );
  XOR2_X2 U5884 ( .A(n3657), .B(n3658), .Z(n3945) );
  XOR2_X2 U5885 ( .A(execstage_BusA[27]), .B(n3656), .Z(n3658) );
  XNOR2_X2 U5886 ( .A(n13132), .B(n16427), .ZN(n3656) );
  OAI22_X2 U5887 ( .A1(n16428), .A2(n8733), .B1(n3950), .B2(n3951), .ZN(n3657)
         );
  AOI221_X2 U5889 ( .B1(n13131), .B2(n3953), .C1(n13218), .C2(
        execstage_BusA[27]), .A(n3426), .ZN(n3793) );
  NAND2_X2 U5890 ( .A1(n3954), .A2(n3955), .ZN(n3426) );
  NAND4_X2 U5892 ( .A1(n3956), .A2(n3957), .A3(n3958), .A4(n3959), .ZN(
        aluout_0[26]) );
  OAI22_X2 U5894 ( .A1(n3962), .A2(n16439), .B1(n16486), .B2(n3964), .ZN(n3961) );
  OAI221_X2 U5898 ( .B1(n13227), .B2(n3811), .C1(n2896), .C2(n8733), .A(n13220), .ZN(n3966) );
  XOR2_X2 U5899 ( .A(n3817), .B(n3816), .Z(n3811) );
  NAND2_X2 U5901 ( .A1(n3818), .A2(n3968), .ZN(n3817) );
  OR3_X2 U5903 ( .A1(n3474), .A2(n13152), .A3(n3969), .ZN(n3818) );
  XNOR2_X2 U5904 ( .A(n3820), .B(n3819), .ZN(n3969) );
  XOR2_X2 U5910 ( .A(n3827), .B(n3825), .Z(n3975) );
  NAND2_X2 U5911 ( .A1(n3826), .A2(n3976), .ZN(n3825) );
  OR3_X2 U5913 ( .A1(n3004), .A2(n13790), .A3(n3977), .ZN(n3826) );
  XNOR2_X2 U5914 ( .A(n3831), .B(n3830), .ZN(n3977) );
  AND3_X2 U5918 ( .A1(n13111), .A2(execstage_BusA[4]), .A3(n3982), .ZN(n3832)
         );
  XOR2_X2 U5919 ( .A(n3836), .B(n3835), .Z(n3982) );
  AND3_X2 U5923 ( .A1(n16406), .A2(n13119), .A3(n3987), .ZN(n3837) );
  XOR2_X2 U5924 ( .A(n3841), .B(n3840), .Z(n3987) );
  NAND2_X2 U5926 ( .A1(n3842), .A2(n3991), .ZN(n3841) );
  OR3_X2 U5928 ( .A1(n3178), .A2(n13154), .A3(n3992), .ZN(n3842) );
  XNOR2_X2 U5929 ( .A(n3846), .B(n3845), .ZN(n3992) );
  NAND2_X2 U5931 ( .A1(n3847), .A2(n3996), .ZN(n3846) );
  OR3_X2 U5933 ( .A1(n3515), .A2(n8739), .A3(n3997), .ZN(n3847) );
  XNOR2_X2 U5934 ( .A(n3851), .B(n3850), .ZN(n3997) );
  NAND2_X2 U5936 ( .A1(n3852), .A2(n4001), .ZN(n3851) );
  OR3_X2 U5938 ( .A1(n3201), .A2(n8714), .A3(n4002), .ZN(n3852) );
  XNOR2_X2 U5939 ( .A(n3856), .B(n3855), .ZN(n4002) );
  NAND2_X2 U5941 ( .A1(n3857), .A2(n4006), .ZN(n3856) );
  OR3_X2 U5943 ( .A1(n3529), .A2(n13146), .A3(n4007), .ZN(n3857) );
  XNOR2_X2 U5944 ( .A(n3861), .B(n3860), .ZN(n4007) );
  NAND2_X2 U5946 ( .A1(n3862), .A2(n4011), .ZN(n3861) );
  OR3_X2 U5948 ( .A1(n13108), .A2(n13136), .A3(n4012), .ZN(n3862) );
  XNOR2_X2 U5949 ( .A(n3866), .B(n3865), .ZN(n4012) );
  NAND2_X2 U5951 ( .A1(n3867), .A2(n4016), .ZN(n3866) );
  OR3_X2 U5953 ( .A1(n3543), .A2(n8736), .A3(n4017), .ZN(n3867) );
  XNOR2_X2 U5954 ( .A(n3872), .B(n3871), .ZN(n4017) );
  NAND2_X2 U5956 ( .A1(n3873), .A2(n4021), .ZN(n3872) );
  OR3_X2 U5958 ( .A1(n13178), .A2(n8695), .A3(n4022), .ZN(n3873) );
  NAND2_X2 U5960 ( .A1(n4023), .A2(n4024), .ZN(n3941) );
  XOR2_X2 U5962 ( .A(n3939), .B(n3940), .Z(n4023) );
  XNOR2_X2 U5963 ( .A(n3879), .B(n3878), .ZN(n3940) );
  NAND2_X2 U5965 ( .A1(n3880), .A2(n4031), .ZN(n3879) );
  OR3_X2 U5967 ( .A1(n8657), .A2(n13162), .A3(n4032), .ZN(n3880) );
  XNOR2_X2 U5968 ( .A(n3884), .B(n3883), .ZN(n4032) );
  AND3_X2 U5973 ( .A1(execstage_BusA[15]), .A2(n13182), .A3(n4038), .ZN(n3885)
         );
  XOR2_X2 U5974 ( .A(n3936), .B(n3937), .Z(n4038) );
  NAND2_X2 U5975 ( .A1(n3938), .A2(n4039), .ZN(n3937) );
  OR3_X2 U5977 ( .A1(n8734), .A2(n13159), .A3(n4040), .ZN(n3938) );
  XNOR2_X2 U5978 ( .A(n3933), .B(n3934), .ZN(n4040) );
  NAND2_X2 U5979 ( .A1(n3935), .A2(n4041), .ZN(n3934) );
  OR3_X2 U5981 ( .A1(n8647), .A2(n13157), .A3(n4042), .ZN(n3935) );
  XNOR2_X2 U5982 ( .A(n3930), .B(n3931), .ZN(n4042) );
  NAND2_X2 U5983 ( .A1(n3932), .A2(n4043), .ZN(n3931) );
  OR3_X2 U5985 ( .A1(n8650), .A2(n13215), .A3(n4044), .ZN(n3932) );
  XNOR2_X2 U5986 ( .A(n3927), .B(n3928), .ZN(n4044) );
  NAND2_X2 U5987 ( .A1(n3929), .A2(n4045), .ZN(n3928) );
  OR3_X2 U5989 ( .A1(n8654), .A2(n13212), .A3(n4046), .ZN(n3929) );
  XNOR2_X2 U5990 ( .A(n3924), .B(n3925), .ZN(n4046) );
  NAND2_X2 U5991 ( .A1(n3926), .A2(n4047), .ZN(n3925) );
  OR3_X2 U5993 ( .A1(n13117), .A2(n13209), .A3(n4048), .ZN(n3926) );
  XNOR2_X2 U5994 ( .A(n3921), .B(n3922), .ZN(n4048) );
  NAND2_X2 U5995 ( .A1(n3923), .A2(n4049), .ZN(n3922) );
  OR3_X2 U5997 ( .A1(n8646), .A2(n13205), .A3(n4050), .ZN(n3923) );
  XOR2_X2 U5998 ( .A(n3920), .B(n3918), .Z(n4050) );
  NAND2_X2 U5999 ( .A1(n3919), .A2(n4051), .ZN(n3918) );
  OR3_X2 U6001 ( .A1(n8653), .A2(n13190), .A3(n4052), .ZN(n3919) );
  XNOR2_X2 U6002 ( .A(n3914), .B(n3915), .ZN(n4052) );
  AND3_X2 U6005 ( .A1(execstage_BusA[23]), .A2(n13204), .A3(n4054), .ZN(n3916)
         );
  XOR2_X2 U6006 ( .A(n3911), .B(n3912), .Z(n4054) );
  NAND2_X2 U6012 ( .A1(n4058), .A2(n4059), .ZN(n3910) );
  XOR2_X2 U6015 ( .A(n3909), .B(n3908), .Z(n4058) );
  NAND2_X2 U6016 ( .A1(execstage_BusA[25]), .A2(n13199), .ZN(n3909) );
  XOR2_X2 U6029 ( .A(n3951), .B(n3950), .Z(n4096) );
  AOI22_X2 U6030 ( .A1(n4097), .A2(execstage_BusA[25]), .B1(n4098), .B2(n4099), 
        .ZN(n3950) );
  XOR2_X2 U6031 ( .A(n8733), .B(n3952), .Z(n3951) );
  XNOR2_X2 U6032 ( .A(n13132), .B(n16429), .ZN(n3952) );
  AOI22_X2 U6035 ( .A1(n16538), .A2(n13196), .B1(execstage_BusA[24]), .B2(
        n13187), .ZN(n4102) );
  NAND4_X2 U6037 ( .A1(n4106), .A2(n4107), .A3(n4108), .A4(n4109), .ZN(
        aluout_0[25]) );
  OAI22_X2 U6039 ( .A1(n16470), .A2(n16439), .B1(n16491), .B2(n3964), .ZN(
        n4111) );
  OAI22_X2 U6042 ( .A1(n16492), .A2(n13103), .B1(n16515), .B2(n2873), .ZN(
        n2706) );
  OAI221_X2 U6045 ( .B1(n13226), .B2(n3967), .C1(n2896), .C2(n8732), .A(n13220), .ZN(n4117) );
  XOR2_X2 U6046 ( .A(n3971), .B(n3970), .Z(n3967) );
  NAND2_X2 U6048 ( .A1(n3972), .A2(n4119), .ZN(n3971) );
  OR3_X2 U6050 ( .A1(n3480), .A2(n13152), .A3(n4120), .ZN(n3972) );
  NAND2_X2 U6052 ( .A1(n4121), .A2(n4122), .ZN(n4094) );
  XOR2_X2 U6054 ( .A(n4093), .B(n4092), .Z(n4121) );
  XNOR2_X2 U6055 ( .A(n3979), .B(n3978), .ZN(n4092) );
  NAND2_X2 U6057 ( .A1(n3980), .A2(n4129), .ZN(n3979) );
  OR3_X2 U6059 ( .A1(n3494), .A2(n13790), .A3(n4130), .ZN(n3980) );
  XNOR2_X2 U6060 ( .A(n3984), .B(n3983), .ZN(n4130) );
  NAND2_X2 U6062 ( .A1(n3985), .A2(n4134), .ZN(n3984) );
  OR3_X2 U6064 ( .A1(n3500), .A2(n8738), .A3(n4135), .ZN(n3985) );
  XNOR2_X2 U6065 ( .A(n3989), .B(n3988), .ZN(n4135) );
  AND3_X2 U6069 ( .A1(n16409), .A2(execstage_BusA[5]), .A3(n4140), .ZN(n3990)
         );
  XOR2_X2 U6070 ( .A(n3994), .B(n3993), .Z(n4140) );
  AND3_X2 U6074 ( .A1(n13112), .A2(n13116), .A3(n4145), .ZN(n3995) );
  XOR2_X2 U6075 ( .A(n3999), .B(n3998), .Z(n4145) );
  AND3_X2 U6079 ( .A1(n13109), .A2(execstage_BusA[7]), .A3(n4150), .ZN(n4000)
         );
  XOR2_X2 U6080 ( .A(n4004), .B(n4003), .Z(n4150) );
  AND3_X2 U6084 ( .A1(n13113), .A2(execstage_BusA[8]), .A3(n4155), .ZN(n4005)
         );
  XOR2_X2 U6085 ( .A(n4009), .B(n4008), .Z(n4155) );
  AND3_X2 U6089 ( .A1(n13107), .A2(n13118), .A3(n4160), .ZN(n4010) );
  XOR2_X2 U6090 ( .A(n4014), .B(n4013), .Z(n4160) );
  AND3_X2 U6094 ( .A1(n13168), .A2(n8694), .A3(n4165), .ZN(n4015) );
  XOR2_X2 U6095 ( .A(n4019), .B(n4018), .Z(n4165) );
  AND3_X2 U6099 ( .A1(n13179), .A2(n13121), .A3(n4170), .ZN(n4020) );
  XOR2_X2 U6100 ( .A(n4026), .B(n16269), .Z(n4170) );
  NAND2_X2 U6103 ( .A1(n4027), .A2(n4175), .ZN(n4026) );
  OR3_X2 U6105 ( .A1(n13165), .A2(n8695), .A3(n4176), .ZN(n4027) );
  XNOR2_X2 U6106 ( .A(n4028), .B(n4029), .ZN(n4176) );
  AND3_X2 U6109 ( .A1(n8655), .A2(n13164), .A3(n4178), .ZN(n4030) );
  XNOR2_X2 U6110 ( .A(n4036), .B(n4034), .ZN(n4178) );
  NAND2_X2 U6111 ( .A1(n4035), .A2(n4179), .ZN(n4034) );
  OR3_X2 U6113 ( .A1(n8657), .A2(n3130), .A3(n4180), .ZN(n4035) );
  XNOR2_X2 U6114 ( .A(n4089), .B(n4090), .ZN(n4180) );
  AND3_X2 U6117 ( .A1(execstage_BusA[15]), .A2(n13161), .A3(n4182), .ZN(n4091)
         );
  XOR2_X2 U6118 ( .A(n4086), .B(n4087), .Z(n4182) );
  AND3_X2 U6121 ( .A1(execstage_BusA[16]), .A2(n13158), .A3(n4184), .ZN(n4088)
         );
  XOR2_X2 U6122 ( .A(n4083), .B(n4084), .Z(n4184) );
  AND3_X2 U6125 ( .A1(execstage_BusA[17]), .A2(n13217), .A3(n4186), .ZN(n4085)
         );
  XOR2_X2 U6126 ( .A(n4080), .B(n4081), .Z(n4186) );
  AND3_X2 U6129 ( .A1(execstage_BusA[18]), .A2(n13214), .A3(n4188), .ZN(n4082)
         );
  XOR2_X2 U6130 ( .A(n4077), .B(n4078), .Z(n4188) );
  AND3_X2 U6133 ( .A1(execstage_BusA[19]), .A2(n13211), .A3(n4190), .ZN(n4079)
         );
  XOR2_X2 U6134 ( .A(n4074), .B(n4075), .Z(n4190) );
  AND3_X2 U6137 ( .A1(execstage_BusA[20]), .A2(n13208), .A3(n4192), .ZN(n4076)
         );
  XNOR2_X2 U6138 ( .A(n4073), .B(n4071), .ZN(n4192) );
  XOR2_X2 U6141 ( .A(n16377), .B(n4068), .Z(n4194) );
  NAND2_X2 U6142 ( .A1(n4069), .A2(n4195), .ZN(n4068) );
  OR3_X2 U6144 ( .A1(n8653), .A2(n13201), .A3(n4196), .ZN(n4069) );
  XNOR2_X2 U6145 ( .A(n4065), .B(n16381), .ZN(n4196) );
  NAND2_X2 U6149 ( .A1(n4066), .A2(n4202), .ZN(n4065) );
  OR3_X2 U6151 ( .A1(n8656), .A2(n13174), .A3(n4203), .ZN(n4066) );
  XOR2_X2 U6152 ( .A(n4063), .B(n4061), .Z(n4203) );
  NAND2_X2 U6153 ( .A1(n4062), .A2(n4204), .ZN(n4061) );
  NAND2_X2 U6155 ( .A1(n3638), .A2(execstage_BusA[24]), .ZN(n4062) );
  NAND2_X2 U6169 ( .A1(n16431), .A2(n13792), .ZN(n4093) );
  OAI221_X2 U6171 ( .B1(n13186), .B2(n8656), .C1(n13170), .C2(n8732), .A(n4240), .ZN(n3440) );
  AOI22_X2 U6172 ( .A1(n16526), .A2(n13198), .B1(n16527), .B2(n13195), .ZN(
        n4240) );
  OAI222_X2 U6173 ( .A1(n16488), .A2(n13104), .B1(n16489), .B2(n2873), .C1(
        n16490), .C2(n13103), .ZN(n2732) );
  OAI221_X2 U6174 ( .B1(n16492), .B2(n13103), .C1(n16517), .C2(n2873), .A(
        n4245), .ZN(n2734) );
  XOR2_X2 U6177 ( .A(n4098), .B(n4099), .Z(n4247) );
  XOR2_X2 U6178 ( .A(execstage_BusA[25]), .B(n4097), .Z(n4099) );
  XNOR2_X2 U6179 ( .A(n13132), .B(n16435), .ZN(n4097) );
  OAI22_X2 U6180 ( .A1(n16432), .A2(n8731), .B1(n4250), .B2(n4251), .ZN(n4098)
         );
  NAND4_X2 U6182 ( .A1(n4253), .A2(n4254), .A3(n4255), .A4(n4256), .ZN(
        aluout_0[24]) );
  OAI22_X2 U6184 ( .A1(n2746), .A2(n4259), .B1(n16493), .B2(n3964), .ZN(n4258)
         );
  AOI22_X2 U6186 ( .A1(n3652), .A2(n16471), .B1(n4261), .B2(n8659), .ZN(n2746)
         );
  OAI221_X2 U6189 ( .B1(n13227), .B2(n4118), .C1(n2896), .C2(n8731), .A(n13220), .ZN(n4263) );
  XOR2_X2 U6190 ( .A(n4124), .B(n4123), .Z(n4118) );
  NAND2_X2 U6192 ( .A1(n4125), .A2(n4265), .ZN(n4124) );
  OR3_X2 U6194 ( .A1(n3004), .A2(n13152), .A3(n4266), .ZN(n4125) );
  XNOR2_X2 U6195 ( .A(n4127), .B(n4126), .ZN(n4266) );
  AND3_X2 U6199 ( .A1(n13111), .A2(n13792), .A3(n4271), .ZN(n4128) );
  XOR2_X2 U6200 ( .A(n4131), .B(n4132), .Z(n4271) );
  AND3_X2 U6203 ( .A1(n16406), .A2(n13791), .A3(n4273), .ZN(n4133) );
  XOR2_X2 U6204 ( .A(n4137), .B(n16198), .Z(n4273) );
  NAND2_X2 U6207 ( .A1(n4138), .A2(n4278), .ZN(n4137) );
  OR3_X2 U6209 ( .A1(n3178), .A2(n8738), .A3(n4279), .ZN(n4138) );
  XNOR2_X2 U6210 ( .A(n4142), .B(n16199), .ZN(n4279) );
  NAND2_X2 U6213 ( .A1(n4143), .A2(n4284), .ZN(n4142) );
  OR3_X2 U6215 ( .A1(n3515), .A2(n13143), .A3(n4285), .ZN(n4143) );
  XNOR2_X2 U6216 ( .A(n4147), .B(n16203), .ZN(n4285) );
  NAND2_X2 U6219 ( .A1(n4148), .A2(n4290), .ZN(n4147) );
  OR3_X2 U6221 ( .A1(n3201), .A2(n13154), .A3(n4291), .ZN(n4148) );
  XNOR2_X2 U6222 ( .A(n4152), .B(n16206), .ZN(n4291) );
  NAND2_X2 U6225 ( .A1(n4153), .A2(n4296), .ZN(n4152) );
  OR3_X2 U6227 ( .A1(n3529), .A2(n13155), .A3(n4297), .ZN(n4153) );
  XNOR2_X2 U6228 ( .A(n4157), .B(n16266), .ZN(n4297) );
  NAND2_X2 U6231 ( .A1(n4158), .A2(n4302), .ZN(n4157) );
  OR3_X2 U6233 ( .A1(n3145), .A2(n13148), .A3(n4303), .ZN(n4158) );
  XNOR2_X2 U6234 ( .A(n4162), .B(n16267), .ZN(n4303) );
  NAND2_X2 U6237 ( .A1(n4163), .A2(n4308), .ZN(n4162) );
  OR3_X2 U6239 ( .A1(n3543), .A2(n13146), .A3(n4309), .ZN(n4163) );
  XNOR2_X2 U6240 ( .A(n4167), .B(n16268), .ZN(n4309) );
  NAND2_X2 U6243 ( .A1(n4168), .A2(n4314), .ZN(n4167) );
  OR3_X2 U6245 ( .A1(n13178), .A2(n13136), .A3(n4315), .ZN(n4168) );
  XNOR2_X2 U6246 ( .A(n4173), .B(n16270), .ZN(n4315) );
  NAND2_X2 U6249 ( .A1(n4174), .A2(n4320), .ZN(n4173) );
  OR3_X2 U6251 ( .A1(n13165), .A2(n8736), .A3(n4321), .ZN(n4174) );
  NAND2_X2 U6253 ( .A1(n4322), .A2(n4323), .ZN(n4239) );
  XOR2_X2 U6255 ( .A(n4237), .B(n4238), .Z(n4322) );
  XNOR2_X2 U6256 ( .A(n4235), .B(n4234), .ZN(n4238) );
  NAND2_X2 U6258 ( .A1(n4236), .A2(n4330), .ZN(n4235) );
  OR3_X2 U6260 ( .A1(n8710), .A2(n3130), .A3(n4331), .ZN(n4236) );
  XNOR2_X2 U6261 ( .A(n4231), .B(n4232), .ZN(n4331) );
  NAND2_X2 U6262 ( .A1(n4233), .A2(n4332), .ZN(n4232) );
  OR3_X2 U6264 ( .A1(n8657), .A2(n13159), .A3(n4333), .ZN(n4233) );
  XNOR2_X2 U6265 ( .A(n4228), .B(n4229), .ZN(n4333) );
  NAND2_X2 U6266 ( .A1(n4230), .A2(n4334), .ZN(n4229) );
  OR3_X2 U6268 ( .A1(n8645), .A2(n13157), .A3(n4335), .ZN(n4230) );
  XNOR2_X2 U6269 ( .A(n4225), .B(n4226), .ZN(n4335) );
  NAND2_X2 U6270 ( .A1(n4227), .A2(n4336), .ZN(n4226) );
  OR3_X2 U6272 ( .A1(n8734), .A2(n13215), .A3(n4337), .ZN(n4227) );
  XNOR2_X2 U6273 ( .A(n4222), .B(n4223), .ZN(n4337) );
  NAND2_X2 U6274 ( .A1(n4224), .A2(n4338), .ZN(n4223) );
  OR3_X2 U6276 ( .A1(n8647), .A2(n13212), .A3(n4339), .ZN(n4224) );
  XNOR2_X2 U6277 ( .A(n4219), .B(n4220), .ZN(n4339) );
  NAND2_X2 U6278 ( .A1(n4221), .A2(n4340), .ZN(n4220) );
  OR3_X2 U6280 ( .A1(n8650), .A2(n13209), .A3(n4341), .ZN(n4221) );
  XNOR2_X2 U6281 ( .A(n4216), .B(n4217), .ZN(n4341) );
  NAND2_X2 U6282 ( .A1(n4218), .A2(n4342), .ZN(n4217) );
  OR3_X2 U6284 ( .A1(n8654), .A2(n13205), .A3(n4343), .ZN(n4218) );
  XNOR2_X2 U6285 ( .A(n4213), .B(n4214), .ZN(n4343) );
  NAND2_X2 U6286 ( .A1(n4215), .A2(n4344), .ZN(n4214) );
  OR3_X2 U6288 ( .A1(n13117), .A2(n13190), .A3(n4345), .ZN(n4215) );
  XNOR2_X2 U6289 ( .A(n4210), .B(n4211), .ZN(n4345) );
  NAND2_X2 U6290 ( .A1(n4212), .A2(n4346), .ZN(n4211) );
  OR3_X2 U6292 ( .A1(n8646), .A2(n13201), .A3(n4347), .ZN(n4212) );
  XOR2_X2 U6293 ( .A(n4201), .B(n4199), .Z(n4347) );
  NAND2_X2 U6294 ( .A1(n4200), .A2(n4348), .ZN(n4199) );
  OR3_X2 U6296 ( .A1(n8653), .A2(n13175), .A3(n4349), .ZN(n4200) );
  NAND2_X2 U6298 ( .A1(n4350), .A2(n4351), .ZN(n4208) );
  XOR2_X2 U6301 ( .A(n4207), .B(n4206), .Z(n4350) );
  NAND2_X2 U6302 ( .A1(execstage_BusA[23]), .A2(n13199), .ZN(n4207) );
  AOI22_X2 U6317 ( .A1(n16534), .A2(n13196), .B1(execstage_BusA[22]), .B2(
        n13187), .ZN(n4391) );
  XOR2_X2 U6319 ( .A(n4251), .B(n4250), .Z(n4393) );
  AOI22_X2 U6320 ( .A1(n4395), .A2(execstage_BusA[23]), .B1(n4396), .B2(n4397), 
        .ZN(n4250) );
  XOR2_X2 U6321 ( .A(n8731), .B(n4252), .Z(n4251) );
  XNOR2_X2 U6322 ( .A(n13133), .B(n16433), .ZN(n4252) );
  NAND4_X2 U6323 ( .A1(n4398), .A2(n4399), .A3(n4400), .A4(n4401), .ZN(
        aluout_0[23]) );
  OAI22_X2 U6325 ( .A1(n16496), .A2(n3964), .B1(n2784), .B2(n4404), .ZN(n4403)
         );
  OAI221_X2 U6329 ( .B1(n13227), .B2(n4264), .C1(n2896), .C2(n8656), .A(n13220), .ZN(n4407) );
  XOR2_X2 U6330 ( .A(n4268), .B(n4267), .Z(n4264) );
  NAND2_X2 U6332 ( .A1(n4269), .A2(n4409), .ZN(n4268) );
  OR3_X2 U6334 ( .A1(n3494), .A2(n13152), .A3(n4410), .ZN(n4269) );
  NAND2_X2 U6336 ( .A1(n4411), .A2(n4412), .ZN(n4385) );
  XOR2_X2 U6338 ( .A(n4384), .B(n4383), .Z(n4411) );
  XNOR2_X2 U6339 ( .A(n4276), .B(n4275), .ZN(n4383) );
  NAND2_X2 U6341 ( .A1(n4277), .A2(n4419), .ZN(n4276) );
  OR3_X2 U6343 ( .A1(n3178), .A2(n13790), .A3(n4420), .ZN(n4277) );
  XNOR2_X2 U6344 ( .A(n4282), .B(n16200), .ZN(n4420) );
  NAND2_X2 U6347 ( .A1(n4283), .A2(n4425), .ZN(n4282) );
  OR3_X2 U6349 ( .A1(n3515), .A2(n8738), .A3(n4426), .ZN(n4283) );
  XNOR2_X2 U6350 ( .A(n4288), .B(n16204), .ZN(n4426) );
  NAND2_X2 U6353 ( .A1(n4289), .A2(n4431), .ZN(n4288) );
  OR3_X2 U6355 ( .A1(n13110), .A2(n13144), .A3(n4432), .ZN(n4289) );
  XNOR2_X2 U6356 ( .A(n4294), .B(n16207), .ZN(n4432) );
  NAND2_X2 U6359 ( .A1(n4295), .A2(n4437), .ZN(n4294) );
  OR3_X2 U6361 ( .A1(n3529), .A2(n13154), .A3(n4438), .ZN(n4295) );
  XNOR2_X2 U6362 ( .A(n4300), .B(n16272), .ZN(n4438) );
  NAND2_X2 U6365 ( .A1(n4301), .A2(n4443), .ZN(n4300) );
  OR3_X2 U6367 ( .A1(n13108), .A2(n13155), .A3(n4444), .ZN(n4301) );
  XNOR2_X2 U6368 ( .A(n4306), .B(n16274), .ZN(n4444) );
  NAND2_X2 U6371 ( .A1(n4307), .A2(n4449), .ZN(n4306) );
  OR3_X2 U6373 ( .A1(n13167), .A2(n13148), .A3(n4450), .ZN(n4307) );
  XNOR2_X2 U6374 ( .A(n4312), .B(n16276), .ZN(n4450) );
  NAND2_X2 U6377 ( .A1(n4313), .A2(n4455), .ZN(n4312) );
  OR3_X2 U6379 ( .A1(n13178), .A2(n13146), .A3(n4456), .ZN(n4313) );
  XNOR2_X2 U6380 ( .A(n4318), .B(n16278), .ZN(n4456) );
  NAND2_X2 U6383 ( .A1(n4319), .A2(n4461), .ZN(n4318) );
  OR3_X2 U6385 ( .A1(n13165), .A2(n13136), .A3(n4462), .ZN(n4319) );
  XNOR2_X2 U6386 ( .A(n4325), .B(n16280), .ZN(n4462) );
  NAND2_X2 U6389 ( .A1(n4326), .A2(n4467), .ZN(n4325) );
  OR3_X2 U6391 ( .A1(n13162), .A2(n8736), .A3(n4468), .ZN(n4326) );
  XNOR2_X2 U6392 ( .A(n4327), .B(n4328), .ZN(n4468) );
  AND3_X2 U6395 ( .A1(execstage_BusA[12]), .A2(n13182), .A3(n4470), .ZN(n4329)
         );
  XOR2_X2 U6396 ( .A(n4380), .B(n4381), .Z(n4470) );
  AND3_X2 U6399 ( .A1(n13120), .A2(n13161), .A3(n4472), .ZN(n4382) );
  XOR2_X2 U6400 ( .A(n4377), .B(n4378), .Z(n4472) );
  AND3_X2 U6403 ( .A1(execstage_BusA[14]), .A2(n13158), .A3(n4474), .ZN(n4379)
         );
  XOR2_X2 U6404 ( .A(n4374), .B(n4375), .Z(n4474) );
  AND3_X2 U6407 ( .A1(execstage_BusA[15]), .A2(n13217), .A3(n4476), .ZN(n4376)
         );
  XOR2_X2 U6408 ( .A(n4371), .B(n4372), .Z(n4476) );
  AND3_X2 U6411 ( .A1(execstage_BusA[16]), .A2(n13214), .A3(n4478), .ZN(n4373)
         );
  XOR2_X2 U6412 ( .A(n4368), .B(n4369), .Z(n4478) );
  AND3_X2 U6415 ( .A1(execstage_BusA[17]), .A2(n13211), .A3(n4480), .ZN(n4370)
         );
  XOR2_X2 U6416 ( .A(n4365), .B(n4366), .Z(n4480) );
  AND3_X2 U6419 ( .A1(execstage_BusA[18]), .A2(n13208), .A3(n4482), .ZN(n4367)
         );
  XOR2_X2 U6420 ( .A(n4362), .B(n4363), .Z(n4482) );
  AND3_X2 U6423 ( .A1(execstage_BusA[19]), .A2(n13188), .A3(n4484), .ZN(n4364)
         );
  XOR2_X2 U6424 ( .A(n4359), .B(n4360), .Z(n4484) );
  AND3_X2 U6427 ( .A1(execstage_BusA[20]), .A2(n13204), .A3(n4486), .ZN(n4361)
         );
  XOR2_X2 U6428 ( .A(n4356), .B(n4357), .Z(n4486) );
  NAND2_X2 U6429 ( .A1(n4358), .A2(n4487), .ZN(n4357) );
  OR3_X2 U6431 ( .A1(n8646), .A2(n13174), .A3(n4488), .ZN(n4358) );
  XOR2_X2 U6432 ( .A(n4355), .B(n4353), .Z(n4488) );
  NAND2_X2 U6433 ( .A1(n4354), .A2(n4489), .ZN(n4353) );
  NAND2_X2 U6435 ( .A1(n16505), .A2(execstage_BusA[22]), .ZN(n4354) );
  NAND2_X2 U6447 ( .A1(n16406), .A2(n13792), .ZN(n4384) );
  AOI221_X2 U6448 ( .B1(n16455), .B2(n2913), .C1(n4114), .C2(n2779), .A(n16443), .ZN(n4399) );
  AOI22_X2 U6450 ( .A1(n2780), .A2(n3806), .B1(n2916), .B2(n13106), .ZN(n4526)
         );
  OAI221_X2 U6451 ( .B1(n13186), .B2(n8646), .C1(n13170), .C2(n8656), .A(n4527), .ZN(n2916) );
  AOI22_X2 U6452 ( .A1(n16526), .A2(n13195), .B1(n16525), .B2(n13200), .ZN(
        n4527) );
  NAND2_X2 U6453 ( .A1(n4529), .A2(n4245), .ZN(n2780) );
  AOI22_X2 U6455 ( .A1(n3803), .A2(n16471), .B1(n4531), .B2(n8659), .ZN(n4529)
         );
  XOR2_X2 U6457 ( .A(n4396), .B(n4397), .Z(n4532) );
  XOR2_X2 U6458 ( .A(execstage_BusA[23]), .B(n4395), .Z(n4397) );
  XNOR2_X2 U6459 ( .A(n13133), .B(n16431), .ZN(n4395) );
  OAI22_X2 U6460 ( .A1(n16410), .A2(n8653), .B1(n4535), .B2(n4536), .ZN(n4396)
         );
  NAND4_X2 U6462 ( .A1(n4538), .A2(n4539), .A3(n4540), .A4(n4541), .ZN(
        aluout_0[22]) );
  OAI22_X2 U6464 ( .A1(n16503), .A2(n3964), .B1(n16513), .B2(n4404), .ZN(n4543) );
  OAI221_X2 U6467 ( .B1(n13227), .B2(n4408), .C1(n2896), .C2(n8653), .A(n13220), .ZN(n4545) );
  XOR2_X2 U6468 ( .A(n4414), .B(n4413), .Z(n4408) );
  NAND2_X2 U6470 ( .A1(n4415), .A2(n4547), .ZN(n4414) );
  OR3_X2 U6472 ( .A1(n3500), .A2(n13152), .A3(n4548), .ZN(n4415) );
  XNOR2_X2 U6473 ( .A(n4417), .B(n4416), .ZN(n4548) );
  XNOR2_X2 U6479 ( .A(n4423), .B(n16202), .ZN(n4554) );
  NAND2_X2 U6482 ( .A1(n4424), .A2(n4559), .ZN(n4423) );
  OR3_X2 U6484 ( .A1(n3515), .A2(n8740), .A3(n4560), .ZN(n4424) );
  XNOR2_X2 U6485 ( .A(n4429), .B(n16205), .ZN(n4560) );
  NAND2_X2 U6488 ( .A1(n4430), .A2(n4565), .ZN(n4429) );
  OR3_X2 U6490 ( .A1(n13110), .A2(n8738), .A3(n4566), .ZN(n4430) );
  XNOR2_X2 U6491 ( .A(n4435), .B(n16208), .ZN(n4566) );
  NAND2_X2 U6494 ( .A1(n4436), .A2(n4571), .ZN(n4435) );
  OR3_X2 U6496 ( .A1(n3529), .A2(n13144), .A3(n4572), .ZN(n4436) );
  XNOR2_X2 U6497 ( .A(n4441), .B(n16273), .ZN(n4572) );
  NAND2_X2 U6500 ( .A1(n4442), .A2(n4577), .ZN(n4441) );
  OR3_X2 U6502 ( .A1(n13108), .A2(n13154), .A3(n4578), .ZN(n4442) );
  XNOR2_X2 U6503 ( .A(n4447), .B(n16275), .ZN(n4578) );
  NAND2_X2 U6506 ( .A1(n4448), .A2(n4583), .ZN(n4447) );
  OR3_X2 U6508 ( .A1(n3543), .A2(n13155), .A3(n4584), .ZN(n4448) );
  XNOR2_X2 U6509 ( .A(n4453), .B(n16277), .ZN(n4584) );
  NAND2_X2 U6512 ( .A1(n4454), .A2(n4589), .ZN(n4453) );
  OR3_X2 U6514 ( .A1(n13178), .A2(n13148), .A3(n4590), .ZN(n4454) );
  XNOR2_X2 U6515 ( .A(n4459), .B(n16279), .ZN(n4590) );
  NAND2_X2 U6518 ( .A1(n4460), .A2(n4595), .ZN(n4459) );
  OR3_X2 U6520 ( .A1(n13165), .A2(n13146), .A3(n4596), .ZN(n4460) );
  XNOR2_X2 U6521 ( .A(n4465), .B(n16281), .ZN(n4596) );
  NAND2_X2 U6524 ( .A1(n4466), .A2(n4601), .ZN(n4465) );
  OR3_X2 U6526 ( .A1(n13162), .A2(n13136), .A3(n4602), .ZN(n4466) );
  NAND2_X2 U6528 ( .A1(n4603), .A2(n4604), .ZN(n4524) );
  XNOR2_X2 U6530 ( .A(n16369), .B(n4523), .ZN(n4603) );
  XNOR2_X2 U6531 ( .A(n4519), .B(n4520), .ZN(n4523) );
  NAND2_X2 U6532 ( .A1(n4521), .A2(n4609), .ZN(n4520) );
  OR3_X2 U6534 ( .A1(n8695), .A2(n13159), .A3(n4610), .ZN(n4521) );
  XNOR2_X2 U6535 ( .A(n4516), .B(n4517), .ZN(n4610) );
  NAND2_X2 U6536 ( .A1(n4518), .A2(n4611), .ZN(n4517) );
  OR3_X2 U6538 ( .A1(n8710), .A2(n13157), .A3(n4612), .ZN(n4518) );
  XNOR2_X2 U6539 ( .A(n4513), .B(n4514), .ZN(n4612) );
  NAND2_X2 U6540 ( .A1(n4515), .A2(n4613), .ZN(n4514) );
  OR3_X2 U6542 ( .A1(n8657), .A2(n13215), .A3(n4614), .ZN(n4515) );
  XNOR2_X2 U6543 ( .A(n4510), .B(n4511), .ZN(n4614) );
  NAND2_X2 U6544 ( .A1(n4512), .A2(n4615), .ZN(n4511) );
  OR3_X2 U6546 ( .A1(n8645), .A2(n13212), .A3(n4616), .ZN(n4512) );
  XNOR2_X2 U6547 ( .A(n4507), .B(n4508), .ZN(n4616) );
  NAND2_X2 U6548 ( .A1(n4509), .A2(n4617), .ZN(n4508) );
  OR3_X2 U6550 ( .A1(n8734), .A2(n13209), .A3(n4618), .ZN(n4509) );
  XNOR2_X2 U6551 ( .A(n4504), .B(n4505), .ZN(n4618) );
  NAND2_X2 U6552 ( .A1(n4506), .A2(n4619), .ZN(n4505) );
  OR3_X2 U6554 ( .A1(n8647), .A2(n13205), .A3(n4620), .ZN(n4506) );
  XNOR2_X2 U6555 ( .A(n4501), .B(n4502), .ZN(n4620) );
  NAND2_X2 U6556 ( .A1(n4503), .A2(n4621), .ZN(n4502) );
  OR3_X2 U6558 ( .A1(n8650), .A2(n13190), .A3(n4622), .ZN(n4503) );
  XNOR2_X2 U6559 ( .A(n4498), .B(n4499), .ZN(n4622) );
  NAND2_X2 U6560 ( .A1(n4500), .A2(n4623), .ZN(n4499) );
  OR3_X2 U6562 ( .A1(n8654), .A2(n13201), .A3(n4624), .ZN(n4500) );
  XNOR2_X2 U6563 ( .A(n4495), .B(n4496), .ZN(n4624) );
  NAND2_X2 U6569 ( .A1(n4628), .A2(n4629), .ZN(n4494) );
  XOR2_X2 U6572 ( .A(n4493), .B(n4492), .Z(n4628) );
  NAND2_X2 U6573 ( .A1(execstage_BusA[21]), .A2(n13199), .ZN(n4493) );
  AOI221_X2 U6583 ( .B1(n13105), .B2(n3237), .C1(n3806), .C2(n2809), .A(n16442), .ZN(n4539) );
  AOI22_X2 U6585 ( .A1(n2808), .A2(n4114), .B1(n3235), .B2(n16455), .ZN(n4662)
         );
  OAI211_X2 U6587 ( .C1(n16519), .C2(n13104), .A(n4666), .B(n4664), .ZN(n2809)
         );
  AOI22_X2 U6588 ( .A1(n4667), .A2(n16471), .B1(n4668), .B2(n8659), .ZN(n4664)
         );
  OAI221_X2 U6589 ( .B1(n13185), .B2(n8730), .C1(n13170), .C2(n8653), .A(n4669), .ZN(n3237) );
  AOI22_X2 U6590 ( .A1(n16404), .A2(n13197), .B1(n16535), .B2(n13195), .ZN(
        n4669) );
  XOR2_X2 U6592 ( .A(n4536), .B(n4535), .Z(n4672) );
  AOI22_X2 U6593 ( .A1(n4674), .A2(execstage_BusA[21]), .B1(n4675), .B2(n4676), 
        .ZN(n4535) );
  XOR2_X2 U6594 ( .A(n8653), .B(n4537), .Z(n4536) );
  XNOR2_X2 U6595 ( .A(n13133), .B(n13111), .ZN(n4537) );
  NAND4_X2 U6596 ( .A1(n4677), .A2(n4678), .A3(n4679), .A4(n4680), .ZN(
        aluout_0[21]) );
  OAI22_X2 U6598 ( .A1(n16490), .A2(n3964), .B1(n16488), .B2(n4404), .ZN(n4682) );
  NAND2_X2 U6599 ( .A1(n16471), .A2(n3808), .ZN(n4404) );
  OAI221_X2 U6602 ( .B1(n13227), .B2(n4546), .C1(n2896), .C2(n8646), .A(n13220), .ZN(n4684) );
  XOR2_X2 U6603 ( .A(n4550), .B(n4549), .Z(n4546) );
  NAND2_X2 U6605 ( .A1(n4551), .A2(n4686), .ZN(n4550) );
  OR3_X2 U6607 ( .A1(n3178), .A2(n13152), .A3(n4687), .ZN(n4551) );
  NAND2_X2 U6609 ( .A1(n4688), .A2(n4689), .ZN(n4558) );
  XOR2_X2 U6611 ( .A(n4557), .B(n4556), .Z(n4688) );
  XNOR2_X2 U6612 ( .A(n4563), .B(n4562), .ZN(n4556) );
  NAND2_X2 U6614 ( .A1(n4564), .A2(n4696), .ZN(n4563) );
  OR3_X2 U6616 ( .A1(n3201), .A2(n13790), .A3(n4697), .ZN(n4564) );
  XNOR2_X2 U6617 ( .A(n4569), .B(n4568), .ZN(n4697) );
  NAND2_X2 U6619 ( .A1(n4570), .A2(n4701), .ZN(n4569) );
  OR3_X2 U6621 ( .A1(n3529), .A2(n8738), .A3(n4702), .ZN(n4570) );
  XNOR2_X2 U6622 ( .A(n4575), .B(n16282), .ZN(n4702) );
  NAND2_X2 U6625 ( .A1(n4576), .A2(n4707), .ZN(n4575) );
  OR3_X2 U6627 ( .A1(n3145), .A2(n13144), .A3(n4708), .ZN(n4576) );
  XNOR2_X2 U6628 ( .A(n4581), .B(n16284), .ZN(n4708) );
  NAND2_X2 U6631 ( .A1(n4582), .A2(n4713), .ZN(n4581) );
  OR3_X2 U6633 ( .A1(n3543), .A2(n13154), .A3(n4714), .ZN(n4582) );
  XNOR2_X2 U6634 ( .A(n4587), .B(n16286), .ZN(n4714) );
  NAND2_X2 U6637 ( .A1(n4588), .A2(n4719), .ZN(n4587) );
  OR3_X2 U6639 ( .A1(n13178), .A2(n13155), .A3(n4720), .ZN(n4588) );
  XNOR2_X2 U6640 ( .A(n4593), .B(n16288), .ZN(n4720) );
  NAND2_X2 U6643 ( .A1(n4594), .A2(n4725), .ZN(n4593) );
  OR3_X2 U6645 ( .A1(n13165), .A2(n13148), .A3(n4726), .ZN(n4594) );
  XNOR2_X2 U6646 ( .A(n4599), .B(n16290), .ZN(n4726) );
  NAND2_X2 U6649 ( .A1(n4600), .A2(n4731), .ZN(n4599) );
  OR3_X2 U6651 ( .A1(n13162), .A2(n13146), .A3(n4732), .ZN(n4600) );
  XNOR2_X2 U6652 ( .A(n4606), .B(n16292), .ZN(n4732) );
  NAND2_X2 U6655 ( .A1(n4607), .A2(n4737), .ZN(n4606) );
  OR3_X2 U6657 ( .A1(n3130), .A2(n13136), .A3(n4738), .ZN(n4607) );
  XNOR2_X2 U6658 ( .A(n4658), .B(n4659), .ZN(n4738) );
  AND3_X2 U6661 ( .A1(n8652), .A2(n13161), .A3(n4740), .ZN(n4660) );
  XOR2_X2 U6662 ( .A(n4655), .B(n4656), .Z(n4740) );
  AND3_X2 U6665 ( .A1(execstage_BusA[12]), .A2(n13158), .A3(n4742), .ZN(n4657)
         );
  XOR2_X2 U6666 ( .A(n4652), .B(n4653), .Z(n4742) );
  AND3_X2 U6669 ( .A1(n8655), .A2(n13217), .A3(n4744), .ZN(n4654) );
  XOR2_X2 U6670 ( .A(n4649), .B(n4650), .Z(n4744) );
  AND3_X2 U6673 ( .A1(execstage_BusA[14]), .A2(n13214), .A3(n4746), .ZN(n4651)
         );
  XOR2_X2 U6674 ( .A(n4646), .B(n4647), .Z(n4746) );
  AND3_X2 U6677 ( .A1(execstage_BusA[15]), .A2(n13211), .A3(n4748), .ZN(n4648)
         );
  XOR2_X2 U6678 ( .A(n4643), .B(n4644), .Z(n4748) );
  AND3_X2 U6681 ( .A1(execstage_BusA[16]), .A2(n13208), .A3(n4750), .ZN(n4645)
         );
  XOR2_X2 U6682 ( .A(n4640), .B(n4641), .Z(n4750) );
  AND3_X2 U6685 ( .A1(execstage_BusA[17]), .A2(n13188), .A3(n4752), .ZN(n4642)
         );
  XOR2_X2 U6686 ( .A(n4637), .B(n4638), .Z(n4752) );
  XNOR2_X2 U6691 ( .A(n4635), .B(n16389), .ZN(n4755) );
  NAND2_X2 U6695 ( .A1(n4636), .A2(n4761), .ZN(n4635) );
  OR3_X2 U6697 ( .A1(n8654), .A2(n13175), .A3(n4762), .ZN(n4636) );
  XOR2_X2 U6698 ( .A(n4633), .B(n4631), .Z(n4762) );
  NAND2_X2 U6699 ( .A1(n4632), .A2(n4763), .ZN(n4631) );
  NAND2_X2 U6701 ( .A1(n16502), .A2(execstage_BusA[20]), .ZN(n4632) );
  NAND2_X2 U6711 ( .A1(n13112), .A2(n13792), .ZN(n4557) );
  AOI221_X2 U6712 ( .B1(n13105), .B2(n3439), .C1(n3806), .C2(n2832), .A(n16441), .ZN(n4678) );
  AOI22_X2 U6714 ( .A1(n2831), .A2(n4114), .B1(n3441), .B2(n16455), .ZN(n4794)
         );
  OAI211_X2 U6716 ( .C1(n16517), .C2(n13104), .A(n4666), .B(n4795), .ZN(n2832)
         );
  AOI22_X2 U6717 ( .A1(n4246), .A2(n16471), .B1(n2727), .B2(n8659), .ZN(n4795)
         );
  OAI221_X2 U6718 ( .B1(n13185), .B2(n8654), .C1(n13170), .C2(n8646), .A(n4796), .ZN(n3439) );
  XOR2_X2 U6721 ( .A(n4675), .B(n4676), .Z(n4798) );
  XOR2_X2 U6722 ( .A(execstage_BusA[21]), .B(n4674), .Z(n4676) );
  XNOR2_X2 U6723 ( .A(n13133), .B(n16406), .ZN(n4674) );
  OAI22_X2 U6724 ( .A1(n16407), .A2(n8730), .B1(n4801), .B2(n4802), .ZN(n4675)
         );
  NAND4_X2 U6726 ( .A1(n4804), .A2(n4805), .A3(n4806), .A4(n4807), .ZN(
        aluout_0[20]) );
  AOI221_X2 U6727 ( .B1(n4685), .B2(n4808), .C1(n16453), .C2(n3645), .A(n4809), 
        .ZN(n4807) );
  NAND2_X2 U6728 ( .A1(n4810), .A2(n3954), .ZN(n4809) );
  OAI221_X2 U6738 ( .B1(n13227), .B2(n4685), .C1(n2896), .C2(n8730), .A(n13220), .ZN(n4811) );
  XOR2_X2 U6739 ( .A(n4691), .B(n4690), .Z(n4685) );
  NAND2_X2 U6741 ( .A1(n4692), .A2(n4816), .ZN(n4691) );
  OR3_X2 U6743 ( .A1(n3515), .A2(n13152), .A3(n4817), .ZN(n4692) );
  XNOR2_X2 U6744 ( .A(n4694), .B(n4693), .ZN(n4817) );
  AND3_X2 U6748 ( .A1(n13109), .A2(n13792), .A3(n4822), .ZN(n4695) );
  XOR2_X2 U6749 ( .A(n4698), .B(n4699), .Z(n4822) );
  AND3_X2 U6752 ( .A1(n13113), .A2(n13791), .A3(n4824), .ZN(n4700) );
  XOR2_X2 U6753 ( .A(n4705), .B(n16283), .Z(n4824) );
  NAND2_X2 U6756 ( .A1(n4706), .A2(n4829), .ZN(n4705) );
  OR3_X2 U6758 ( .A1(n13108), .A2(n8738), .A3(n4830), .ZN(n4706) );
  XNOR2_X2 U6759 ( .A(n4711), .B(n16285), .ZN(n4830) );
  NAND2_X2 U6762 ( .A1(n4712), .A2(n4835), .ZN(n4711) );
  OR3_X2 U6764 ( .A1(n3543), .A2(n13144), .A3(n4836), .ZN(n4712) );
  XNOR2_X2 U6765 ( .A(n4717), .B(n16287), .ZN(n4836) );
  NAND2_X2 U6768 ( .A1(n4718), .A2(n4841), .ZN(n4717) );
  OR3_X2 U6770 ( .A1(n13178), .A2(n13154), .A3(n4842), .ZN(n4718) );
  XNOR2_X2 U6771 ( .A(n4723), .B(n16289), .ZN(n4842) );
  NAND2_X2 U6774 ( .A1(n4724), .A2(n4847), .ZN(n4723) );
  OR3_X2 U6776 ( .A1(n13165), .A2(n13155), .A3(n4848), .ZN(n4724) );
  XNOR2_X2 U6777 ( .A(n4729), .B(n16291), .ZN(n4848) );
  NAND2_X2 U6780 ( .A1(n4730), .A2(n4853), .ZN(n4729) );
  OR3_X2 U6782 ( .A1(n13162), .A2(n13148), .A3(n4854), .ZN(n4730) );
  XNOR2_X2 U6783 ( .A(n4735), .B(n16293), .ZN(n4854) );
  NAND2_X2 U6786 ( .A1(n4736), .A2(n4859), .ZN(n4735) );
  OR3_X2 U6788 ( .A1(n3130), .A2(n13146), .A3(n4860), .ZN(n4736) );
  NAND2_X2 U6790 ( .A1(n4861), .A2(n4862), .ZN(n4792) );
  XOR2_X2 U6792 ( .A(n4790), .B(n4791), .Z(n4861) );
  XNOR2_X2 U6793 ( .A(n4787), .B(n4788), .ZN(n4791) );
  NAND2_X2 U6794 ( .A1(n4789), .A2(n4866), .ZN(n4788) );
  OR3_X2 U6796 ( .A1(n8736), .A2(n13157), .A3(n4867), .ZN(n4789) );
  XNOR2_X2 U6797 ( .A(n4784), .B(n4785), .ZN(n4867) );
  NAND2_X2 U6798 ( .A1(n4786), .A2(n4868), .ZN(n4785) );
  OR3_X2 U6800 ( .A1(n8695), .A2(n13215), .A3(n4869), .ZN(n4786) );
  XNOR2_X2 U6801 ( .A(n4781), .B(n4782), .ZN(n4869) );
  NAND2_X2 U6802 ( .A1(n4783), .A2(n4870), .ZN(n4782) );
  OR3_X2 U6804 ( .A1(n8710), .A2(n13212), .A3(n4871), .ZN(n4783) );
  XNOR2_X2 U6805 ( .A(n4778), .B(n4779), .ZN(n4871) );
  NAND2_X2 U6806 ( .A1(n4780), .A2(n4872), .ZN(n4779) );
  OR3_X2 U6808 ( .A1(n8657), .A2(n13209), .A3(n4873), .ZN(n4780) );
  XNOR2_X2 U6809 ( .A(n4775), .B(n4776), .ZN(n4873) );
  NAND2_X2 U6810 ( .A1(n4777), .A2(n4874), .ZN(n4776) );
  OR3_X2 U6812 ( .A1(n8645), .A2(n13205), .A3(n4875), .ZN(n4777) );
  XNOR2_X2 U6813 ( .A(n4772), .B(n4773), .ZN(n4875) );
  NAND2_X2 U6814 ( .A1(n4774), .A2(n4876), .ZN(n4773) );
  OR3_X2 U6816 ( .A1(n8734), .A2(n13190), .A3(n4877), .ZN(n4774) );
  XNOR2_X2 U6817 ( .A(n4769), .B(n4770), .ZN(n4877) );
  NAND2_X2 U6818 ( .A1(n4771), .A2(n4878), .ZN(n4770) );
  OR3_X2 U6820 ( .A1(n8647), .A2(n13201), .A3(n4879), .ZN(n4771) );
  XOR2_X2 U6821 ( .A(n4760), .B(n4758), .Z(n4879) );
  NAND2_X2 U6822 ( .A1(n4759), .A2(n4880), .ZN(n4758) );
  OR3_X2 U6824 ( .A1(n8650), .A2(n13174), .A3(n4881), .ZN(n4759) );
  NAND2_X2 U6826 ( .A1(n4882), .A2(n4883), .ZN(n4768) );
  XOR2_X2 U6828 ( .A(n4767), .B(n4766), .Z(n4882) );
  NAND2_X2 U6829 ( .A1(execstage_BusA[19]), .A2(n13199), .ZN(n4767) );
  OAI221_X2 U6840 ( .B1(n13185), .B2(n8650), .C1(n13170), .C2(n13117), .A(
        n4914), .ZN(n3648) );
  AOI22_X2 U6841 ( .A1(n16404), .A2(n13196), .B1(n16536), .B2(n13200), .ZN(
        n4914) );
  XOR2_X2 U6843 ( .A(n4802), .B(n4801), .Z(n4916) );
  AOI22_X2 U6844 ( .A1(n4918), .A2(execstage_BusA[19]), .B1(n4919), .B2(n4920), 
        .ZN(n4801) );
  XOR2_X2 U6845 ( .A(n8730), .B(n4803), .Z(n4802) );
  XNOR2_X2 U6846 ( .A(n13133), .B(n16409), .ZN(n4803) );
  NAND4_X2 U6847 ( .A1(n4921), .A2(n4922), .A3(n4923), .A4(n4924), .ZN(
        aluout_0[1]) );
  OAI22_X2 U6850 ( .A1(n2827), .A2(n4929), .B1(n4930), .B2(n2772), .ZN(n4926)
         );
  AOI221_X2 U6851 ( .B1(n4931), .B2(n13194), .C1(n13187), .C2(n8651), .A(n4932), .ZN(n4930) );
  AOI221_X2 U6853 ( .B1(execstage_BusA[7]), .B2(n13183), .C1(execstage_BusA[5]), .C2(n13171), .A(n4934), .ZN(n2827) );
  OAI22_X2 U6854 ( .A1(n2885), .A2(n13196), .B1(n2882), .B2(n13200), .ZN(n4934) );
  OAI221_X2 U6856 ( .B1(n13141), .B2(n13185), .C1(n13146), .C2(n13170), .A(
        n4936), .ZN(n2719) );
  AOI22_X2 U6857 ( .A1(n16522), .A2(n13197), .B1(n16529), .B2(n13195), .ZN(
        n4936) );
  XOR2_X2 U6858 ( .A(n4939), .B(n4940), .Z(n4935) );
  AOI221_X2 U6859 ( .B1(n13106), .B2(n4941), .C1(n13223), .C2(n4928), .A(
        n16398), .ZN(n4922) );
  AOI22_X2 U6861 ( .A1(n4944), .A2(n2733), .B1(n4945), .B2(n13114), .ZN(n4943)
         );
  NAND4_X2 U6863 ( .A1(n4949), .A2(n4950), .A3(n4951), .A4(n4952), .ZN(
        aluout_0[19]) );
  OAI22_X2 U6865 ( .A1(n2784), .A2(n4955), .B1(n16495), .B2(n3964), .ZN(n4954)
         );
  OAI221_X2 U6868 ( .B1(n13227), .B2(n4815), .C1(n2896), .C2(n8654), .A(n13220), .ZN(n4956) );
  XOR2_X2 U6869 ( .A(n4819), .B(n4818), .Z(n4815) );
  NAND2_X2 U6871 ( .A1(n4820), .A2(n4958), .ZN(n4819) );
  OR3_X2 U6873 ( .A1(n3201), .A2(n13151), .A3(n4959), .ZN(n4820) );
  NAND2_X2 U6875 ( .A1(n4960), .A2(n4961), .ZN(n4913) );
  XOR2_X2 U6877 ( .A(n4912), .B(n4911), .Z(n4960) );
  XNOR2_X2 U6878 ( .A(n4827), .B(n4826), .ZN(n4911) );
  NAND2_X2 U6880 ( .A1(n4828), .A2(n4968), .ZN(n4827) );
  OR3_X2 U6882 ( .A1(n3145), .A2(n13790), .A3(n4969), .ZN(n4828) );
  XNOR2_X2 U6883 ( .A(n4833), .B(n4832), .ZN(n4969) );
  NAND2_X2 U6885 ( .A1(n4834), .A2(n4973), .ZN(n4833) );
  OR3_X2 U6887 ( .A1(n3543), .A2(n8738), .A3(n4974), .ZN(n4834) );
  XNOR2_X2 U6888 ( .A(n4839), .B(n16297), .ZN(n4974) );
  NAND2_X2 U6891 ( .A1(n4840), .A2(n4979), .ZN(n4839) );
  OR3_X2 U6893 ( .A1(n13178), .A2(n13144), .A3(n4980), .ZN(n4840) );
  XNOR2_X2 U6894 ( .A(n4845), .B(n16299), .ZN(n4980) );
  NAND2_X2 U6897 ( .A1(n4846), .A2(n4985), .ZN(n4845) );
  OR3_X2 U6899 ( .A1(n13165), .A2(n13154), .A3(n4986), .ZN(n4846) );
  XNOR2_X2 U6900 ( .A(n4851), .B(n16303), .ZN(n4986) );
  NAND2_X2 U6903 ( .A1(n4852), .A2(n4991), .ZN(n4851) );
  OR3_X2 U6905 ( .A1(n13162), .A2(n13155), .A3(n4992), .ZN(n4852) );
  XNOR2_X2 U6906 ( .A(n4857), .B(n16305), .ZN(n4992) );
  NAND2_X2 U6909 ( .A1(n4858), .A2(n4997), .ZN(n4857) );
  OR3_X2 U6911 ( .A1(n3130), .A2(n13148), .A3(n4998), .ZN(n4858) );
  XNOR2_X2 U6912 ( .A(n4864), .B(n16307), .ZN(n4998) );
  NAND2_X2 U6915 ( .A1(n4865), .A2(n5003), .ZN(n4864) );
  OR3_X2 U6917 ( .A1(n13159), .A2(n13146), .A3(n5004), .ZN(n4865) );
  XNOR2_X2 U6918 ( .A(n4908), .B(n4909), .ZN(n5004) );
  AND3_X2 U6921 ( .A1(n13122), .A2(n13158), .A3(n5006), .ZN(n4910) );
  XOR2_X2 U6922 ( .A(n4905), .B(n4906), .Z(n5006) );
  AND3_X2 U6925 ( .A1(n8652), .A2(n13217), .A3(n5008), .ZN(n4907) );
  XOR2_X2 U6926 ( .A(n4902), .B(n4903), .Z(n5008) );
  AND3_X2 U6929 ( .A1(execstage_BusA[12]), .A2(n13214), .A3(n5010), .ZN(n4904)
         );
  XOR2_X2 U6930 ( .A(n4899), .B(n4900), .Z(n5010) );
  AND3_X2 U6933 ( .A1(n8655), .A2(n13211), .A3(n5012), .ZN(n4901) );
  XOR2_X2 U6934 ( .A(n4896), .B(n4897), .Z(n5012) );
  AND3_X2 U6937 ( .A1(execstage_BusA[14]), .A2(n13207), .A3(n5014), .ZN(n4898)
         );
  XOR2_X2 U6938 ( .A(n4893), .B(n4894), .Z(n5014) );
  AND3_X2 U6941 ( .A1(execstage_BusA[15]), .A2(n13188), .A3(n5016), .ZN(n4895)
         );
  XOR2_X2 U6942 ( .A(n4890), .B(n4891), .Z(n5016) );
  AND3_X2 U6945 ( .A1(execstage_BusA[16]), .A2(n13204), .A3(n5018), .ZN(n4892)
         );
  XOR2_X2 U6946 ( .A(n4887), .B(n4888), .Z(n5018) );
  NAND2_X2 U6947 ( .A1(n4889), .A2(n5019), .ZN(n4888) );
  OR3_X2 U6949 ( .A1(n8647), .A2(n13174), .A3(n5020), .ZN(n4889) );
  NAND2_X2 U6951 ( .A1(n5021), .A2(n5022), .ZN(n4886) );
  XOR2_X2 U6954 ( .A(n4885), .B(n4884), .Z(n5021) );
  NAND2_X2 U6955 ( .A1(execstage_BusA[18]), .A2(n13198), .ZN(n4885) );
  NAND2_X2 U6964 ( .A1(n13113), .A2(n13792), .ZN(n4912) );
  OAI221_X2 U6966 ( .B1(n13185), .B2(n8647), .C1(n13169), .C2(n8654), .A(
        n16482), .ZN(n2913) );
  OAI211_X2 U6970 ( .C1(n16494), .C2(n13104), .A(n4666), .B(n5055), .ZN(n2893)
         );
  AOI22_X2 U6971 ( .A1(n4531), .A2(n16471), .B1(n2776), .B2(n8659), .ZN(n5055)
         );
  NAND2_X2 U6972 ( .A1(n16469), .A2(execstage_ALU_ra_row2_31_), .ZN(n4666) );
  XOR2_X2 U6974 ( .A(n4919), .B(n4920), .Z(n5057) );
  XOR2_X2 U6975 ( .A(execstage_BusA[19]), .B(n4918), .Z(n4920) );
  XNOR2_X2 U6976 ( .A(n13133), .B(n13112), .ZN(n4918) );
  OAI22_X2 U6977 ( .A1(n16412), .A2(n8650), .B1(n5060), .B2(n5061), .ZN(n4919)
         );
  NAND4_X2 U6979 ( .A1(n5063), .A2(n5064), .A3(n5065), .A4(n5066), .ZN(
        aluout_0[18]) );
  OAI22_X2 U6981 ( .A1(n16513), .A2(n4955), .B1(n16514), .B2(n3964), .ZN(n5068) );
  OAI221_X2 U6984 ( .B1(n13227), .B2(n4957), .C1(n2896), .C2(n8650), .A(n13220), .ZN(n5070) );
  XOR2_X2 U6985 ( .A(n4963), .B(n4962), .Z(n4957) );
  NAND2_X2 U6987 ( .A1(n4964), .A2(n5073), .ZN(n4963) );
  OR3_X2 U6989 ( .A1(n3529), .A2(n13151), .A3(n5074), .ZN(n4964) );
  XNOR2_X2 U6990 ( .A(n4966), .B(n4965), .ZN(n5074) );
  AND3_X2 U6994 ( .A1(n13107), .A2(n13792), .A3(n5079), .ZN(n4967) );
  XOR2_X2 U6995 ( .A(n4970), .B(n4971), .Z(n5079) );
  AND3_X2 U6998 ( .A1(n13168), .A2(n13791), .A3(n5081), .ZN(n4972) );
  XOR2_X2 U6999 ( .A(n4977), .B(n4976), .Z(n5081) );
  NAND2_X2 U7001 ( .A1(n4978), .A2(n5085), .ZN(n4977) );
  OR3_X2 U7003 ( .A1(n13178), .A2(n8738), .A3(n5086), .ZN(n4978) );
  XNOR2_X2 U7004 ( .A(n4983), .B(n16300), .ZN(n5086) );
  NAND2_X2 U7007 ( .A1(n4984), .A2(n5091), .ZN(n4983) );
  OR3_X2 U7009 ( .A1(n13165), .A2(n13144), .A3(n5092), .ZN(n4984) );
  XNOR2_X2 U7010 ( .A(n4989), .B(n16304), .ZN(n5092) );
  NAND2_X2 U7013 ( .A1(n4990), .A2(n5097), .ZN(n4989) );
  OR3_X2 U7015 ( .A1(n13162), .A2(n13154), .A3(n5098), .ZN(n4990) );
  XNOR2_X2 U7016 ( .A(n4995), .B(n16306), .ZN(n5098) );
  NAND2_X2 U7019 ( .A1(n4996), .A2(n5103), .ZN(n4995) );
  OR3_X2 U7021 ( .A1(n3130), .A2(n13155), .A3(n5104), .ZN(n4996) );
  XNOR2_X2 U7022 ( .A(n5001), .B(n16308), .ZN(n5104) );
  NAND2_X2 U7025 ( .A1(n5002), .A2(n5109), .ZN(n5001) );
  OR3_X2 U7027 ( .A1(n13159), .A2(n13148), .A3(n5110), .ZN(n5002) );
  NAND2_X2 U7029 ( .A1(n5111), .A2(n5112), .ZN(n5050) );
  XOR2_X2 U7031 ( .A(n5048), .B(n5049), .Z(n5111) );
  XNOR2_X2 U7032 ( .A(n5045), .B(n5046), .ZN(n5049) );
  NAND2_X2 U7033 ( .A1(n5047), .A2(n5116), .ZN(n5046) );
  OR3_X2 U7035 ( .A1(n13136), .A2(n13215), .A3(n5117), .ZN(n5047) );
  XNOR2_X2 U7036 ( .A(n5042), .B(n5043), .ZN(n5117) );
  NAND2_X2 U7037 ( .A1(n5044), .A2(n5118), .ZN(n5043) );
  OR3_X2 U7039 ( .A1(n8736), .A2(n13212), .A3(n5119), .ZN(n5044) );
  XNOR2_X2 U7040 ( .A(n5039), .B(n5040), .ZN(n5119) );
  NAND2_X2 U7041 ( .A1(n5041), .A2(n5120), .ZN(n5040) );
  OR3_X2 U7043 ( .A1(n8695), .A2(n13209), .A3(n5121), .ZN(n5041) );
  XNOR2_X2 U7044 ( .A(n5036), .B(n5037), .ZN(n5121) );
  NAND2_X2 U7045 ( .A1(n5038), .A2(n5122), .ZN(n5037) );
  OR3_X2 U7047 ( .A1(n8710), .A2(n13205), .A3(n5123), .ZN(n5038) );
  XNOR2_X2 U7048 ( .A(n5033), .B(n5034), .ZN(n5123) );
  NAND2_X2 U7049 ( .A1(n5035), .A2(n5124), .ZN(n5034) );
  OR3_X2 U7051 ( .A1(n8657), .A2(n2909), .A3(n5125), .ZN(n5035) );
  XNOR2_X2 U7052 ( .A(n5030), .B(n5031), .ZN(n5125) );
  NAND2_X2 U7053 ( .A1(n5032), .A2(n5126), .ZN(n5031) );
  OR3_X2 U7055 ( .A1(n8645), .A2(n13201), .A3(n5127), .ZN(n5032) );
  XNOR2_X2 U7056 ( .A(n5027), .B(n5028), .ZN(n5127) );
  AND3_X2 U7059 ( .A1(execstage_BusA[16]), .A2(n13177), .A3(n5129), .ZN(n5029)
         );
  XNOR2_X2 U7060 ( .A(n5026), .B(n5024), .ZN(n5129) );
  NAND2_X2 U7061 ( .A1(n5025), .A2(n5130), .ZN(n5024) );
  NAND2_X2 U7063 ( .A1(n4797), .A2(execstage_BusA[17]), .ZN(n5025) );
  OAI221_X2 U7074 ( .B1(n13139), .B2(n13185), .C1(n13169), .C2(n8650), .A(
        n5158), .ZN(n3235) );
  AOI22_X2 U7075 ( .A1(n16544), .A2(n13197), .B1(n16536), .B2(n13195), .ZN(
        n5158) );
  XOR2_X2 U7081 ( .A(n5061), .B(n5060), .Z(n5162) );
  AOI22_X2 U7082 ( .A1(n5164), .A2(execstage_BusA[17]), .B1(n5165), .B2(n5166), 
        .ZN(n5060) );
  XOR2_X2 U7083 ( .A(n8650), .B(n5062), .Z(n5061) );
  XNOR2_X2 U7084 ( .A(n13133), .B(n13109), .ZN(n5062) );
  NAND4_X2 U7086 ( .A1(n5167), .A2(n5168), .A3(n5169), .A4(n5170), .ZN(
        aluout_0[17]) );
  OAI22_X2 U7088 ( .A1(n16488), .A2(n4955), .B1(n16489), .B2(n3964), .ZN(n5172) );
  OAI221_X2 U7093 ( .B1(n13227), .B2(n5072), .C1(n2896), .C2(n8647), .A(n13220), .ZN(n5173) );
  XOR2_X2 U7094 ( .A(n5076), .B(n5075), .Z(n5072) );
  NAND2_X2 U7096 ( .A1(n5077), .A2(n5176), .ZN(n5076) );
  OR3_X2 U7098 ( .A1(n3145), .A2(n13151), .A3(n5177), .ZN(n5077) );
  NAND2_X2 U7100 ( .A1(n5178), .A2(n5179), .ZN(n5157) );
  XOR2_X2 U7102 ( .A(n5156), .B(n5155), .Z(n5178) );
  XNOR2_X2 U7103 ( .A(n5083), .B(n5082), .ZN(n5155) );
  AND3_X2 U7107 ( .A1(n13179), .A2(n13791), .A3(n5187), .ZN(n5084) );
  XOR2_X2 U7108 ( .A(n5089), .B(n16301), .Z(n5187) );
  NAND2_X2 U7112 ( .A1(n5090), .A2(n5193), .ZN(n5089) );
  OR3_X2 U7114 ( .A1(n13165), .A2(n8738), .A3(n5194), .ZN(n5090) );
  XNOR2_X2 U7115 ( .A(n5095), .B(n5094), .ZN(n5194) );
  NAND2_X2 U7117 ( .A1(n5096), .A2(n5198), .ZN(n5095) );
  OR3_X2 U7119 ( .A1(n13162), .A2(n13144), .A3(n5199), .ZN(n5096) );
  XNOR2_X2 U7120 ( .A(n5101), .B(n5100), .ZN(n5199) );
  NAND2_X2 U7122 ( .A1(n5102), .A2(n5203), .ZN(n5101) );
  OR3_X2 U7124 ( .A1(n3130), .A2(n13154), .A3(n5204), .ZN(n5102) );
  XNOR2_X2 U7125 ( .A(n5107), .B(n16309), .ZN(n5204) );
  NAND2_X2 U7128 ( .A1(n5108), .A2(n5209), .ZN(n5107) );
  OR3_X2 U7130 ( .A1(n13159), .A2(n13155), .A3(n5210), .ZN(n5108) );
  XNOR2_X2 U7131 ( .A(n5114), .B(n16310), .ZN(n5210) );
  NAND2_X2 U7134 ( .A1(n5115), .A2(n5215), .ZN(n5114) );
  OR3_X2 U7136 ( .A1(n13157), .A2(n8714), .A3(n5216), .ZN(n5115) );
  XNOR2_X2 U7137 ( .A(n5152), .B(n5153), .ZN(n5216) );
  AND3_X2 U7140 ( .A1(n13118), .A2(n13217), .A3(n5218), .ZN(n5154) );
  XOR2_X2 U7141 ( .A(n5149), .B(n5150), .Z(n5218) );
  AND3_X2 U7144 ( .A1(n13122), .A2(n13214), .A3(n5220), .ZN(n5151) );
  XOR2_X2 U7145 ( .A(n5146), .B(n5147), .Z(n5220) );
  AND3_X2 U7148 ( .A1(n8652), .A2(n13211), .A3(n5222), .ZN(n5148) );
  XOR2_X2 U7149 ( .A(n5143), .B(n5144), .Z(n5222) );
  AND3_X2 U7152 ( .A1(execstage_BusA[12]), .A2(n13207), .A3(n5224), .ZN(n5145)
         );
  XOR2_X2 U7153 ( .A(n5140), .B(n5141), .Z(n5224) );
  AND3_X2 U7156 ( .A1(n8655), .A2(n13188), .A3(n5226), .ZN(n5142) );
  XOR2_X2 U7157 ( .A(n5137), .B(n5138), .Z(n5226) );
  XNOR2_X2 U7162 ( .A(n5135), .B(n16473), .ZN(n5229) );
  NAND2_X2 U7165 ( .A1(n5136), .A2(n5234), .ZN(n5135) );
  OR3_X2 U7167 ( .A1(n8645), .A2(n13175), .A3(n5235), .ZN(n5136) );
  NAND2_X2 U7169 ( .A1(n5236), .A2(n16485), .ZN(n5133) );
  AOI22_X2 U7171 ( .A1(n5239), .A2(n5240), .B1(n5241), .B2(n5242), .ZN(n5238)
         );
  XOR2_X2 U7172 ( .A(n5132), .B(n5131), .Z(n5236) );
  NAND2_X2 U7173 ( .A1(execstage_BusA[16]), .A2(n13198), .ZN(n5132) );
  NAND2_X2 U7180 ( .A1(n13168), .A2(n13792), .ZN(n5156) );
  AOI22_X2 U7183 ( .A1(n5240), .A2(n5264), .B1(n16523), .B2(n13200), .ZN(n5263) );
  XOR2_X2 U7191 ( .A(n5165), .B(n5166), .Z(n5267) );
  XOR2_X2 U7192 ( .A(execstage_BusA[17]), .B(n5164), .Z(n5166) );
  XNOR2_X2 U7193 ( .A(n13133), .B(n13113), .ZN(n5164) );
  OAI22_X2 U7194 ( .A1(n16418), .A2(n8734), .B1(n5270), .B2(n5271), .ZN(n5165)
         );
  NAND4_X2 U7196 ( .A1(n5273), .A2(n5274), .A3(n5275), .A4(n5276), .ZN(
        aluout_0[16]) );
  AOI221_X2 U7197 ( .B1(n16453), .B2(n4387), .C1(n5175), .C2(n5277), .A(n16458), .ZN(n5276) );
  OAI221_X2 U7202 ( .B1(n5175), .B2(n13226), .C1(n8734), .C2(n2896), .A(n13220), .ZN(n5278) );
  XOR2_X2 U7203 ( .A(n5181), .B(n5180), .Z(n5175) );
  NAND2_X2 U7205 ( .A1(n5182), .A2(n5280), .ZN(n5181) );
  OR3_X2 U7207 ( .A1(n3543), .A2(n13151), .A3(n5281), .ZN(n5182) );
  XNOR2_X2 U7208 ( .A(n5184), .B(n5183), .ZN(n5281) );
  NAND2_X2 U7210 ( .A1(n5185), .A2(n5285), .ZN(n5184) );
  OR3_X2 U7212 ( .A1(n13178), .A2(n13793), .A3(n5286), .ZN(n5185) );
  XOR2_X2 U7213 ( .A(n5192), .B(n5190), .Z(n5286) );
  NAND2_X2 U7214 ( .A1(n5191), .A2(n5287), .ZN(n5190) );
  OR3_X2 U7216 ( .A1(n13165), .A2(n13790), .A3(n5288), .ZN(n5191) );
  XNOR2_X2 U7217 ( .A(n5196), .B(n5195), .ZN(n5288) );
  AND3_X2 U7221 ( .A1(n13164), .A2(execstage_BusA[4]), .A3(n5293), .ZN(n5197)
         );
  XOR2_X2 U7222 ( .A(n5201), .B(n5200), .Z(n5293) );
  AND3_X2 U7226 ( .A1(n13182), .A2(execstage_BusA[5]), .A3(n5298), .ZN(n5202)
         );
  XOR2_X2 U7227 ( .A(n5207), .B(n5206), .Z(n5298) );
  NAND2_X2 U7229 ( .A1(n5208), .A2(n5302), .ZN(n5207) );
  OR3_X2 U7231 ( .A1(n13159), .A2(n8715), .A3(n5303), .ZN(n5208) );
  XNOR2_X2 U7232 ( .A(n5213), .B(n5212), .ZN(n5303) );
  NAND2_X2 U7234 ( .A1(n5214), .A2(n5307), .ZN(n5213) );
  OR3_X2 U7236 ( .A1(n13157), .A2(n13155), .A3(n5308), .ZN(n5214) );
  NAND2_X2 U7238 ( .A1(n5309), .A2(n5310), .ZN(n5260) );
  XOR2_X2 U7240 ( .A(n5259), .B(n5258), .Z(n5309) );
  XNOR2_X2 U7241 ( .A(n16338), .B(n5256), .ZN(n5258) );
  NAND2_X2 U7242 ( .A1(n5257), .A2(n5314), .ZN(n5256) );
  OR3_X2 U7244 ( .A1(n13146), .A2(n13212), .A3(n5315), .ZN(n5257) );
  XNOR2_X2 U7245 ( .A(n5252), .B(n5253), .ZN(n5315) );
  NAND2_X2 U7246 ( .A1(n5254), .A2(n5316), .ZN(n5253) );
  OR3_X2 U7248 ( .A1(n13136), .A2(n13209), .A3(n5317), .ZN(n5254) );
  XNOR2_X2 U7249 ( .A(n5249), .B(n5250), .ZN(n5317) );
  NAND2_X2 U7250 ( .A1(n5251), .A2(n5318), .ZN(n5250) );
  OR3_X2 U7252 ( .A1(n8736), .A2(n13205), .A3(n5319), .ZN(n5251) );
  XNOR2_X2 U7253 ( .A(n5246), .B(n5247), .ZN(n5319) );
  NAND2_X2 U7254 ( .A1(n5248), .A2(n5320), .ZN(n5247) );
  OR3_X2 U7256 ( .A1(n8695), .A2(n2909), .A3(n5321), .ZN(n5248) );
  XNOR2_X2 U7257 ( .A(n5243), .B(n5244), .ZN(n5321) );
  NAND2_X2 U7258 ( .A1(n5245), .A2(n5322), .ZN(n5244) );
  OR3_X2 U7260 ( .A1(n8710), .A2(n13201), .A3(n5323), .ZN(n5245) );
  XNOR2_X2 U7261 ( .A(n5231), .B(n5232), .ZN(n5323) );
  NAND2_X2 U7262 ( .A1(n5233), .A2(n5324), .ZN(n5232) );
  OR3_X2 U7264 ( .A1(n8657), .A2(n13174), .A3(n5325), .ZN(n5233) );
  XNOR2_X2 U7265 ( .A(n5241), .B(n5242), .ZN(n5325) );
  XOR2_X2 U7266 ( .A(n5240), .B(n5239), .Z(n5242) );
  NAND2_X2 U7278 ( .A1(n8659), .A2(n3808), .ZN(n4955) );
  OAI221_X2 U7281 ( .B1(n13138), .B2(n13185), .C1(n8734), .C2(n3434), .A(n5353), .ZN(n3646) );
  AOI22_X2 U7282 ( .A1(n16544), .A2(n13196), .B1(n16543), .B2(n13197), .ZN(
        n5353) );
  XOR2_X2 U7283 ( .A(n5271), .B(n5270), .Z(n5352) );
  AOI22_X2 U7284 ( .A1(n5355), .A2(execstage_BusA[15]), .B1(n5356), .B2(n5357), 
        .ZN(n5270) );
  XOR2_X2 U7285 ( .A(n13139), .B(n5272), .Z(n5271) );
  XNOR2_X2 U7286 ( .A(n13133), .B(n13107), .ZN(n5272) );
  NAND4_X2 U7288 ( .A1(n5361), .A2(n5362), .A3(n5363), .A4(n5364), .ZN(
        aluout_0[15]) );
  AOI22_X2 U7292 ( .A1(n5368), .A2(n16518), .B1(n5369), .B2(n5279), .ZN(n5367)
         );
  XOR2_X2 U7293 ( .A(n5283), .B(n5282), .Z(n5279) );
  NAND2_X2 U7300 ( .A1(n5375), .A2(n5376), .ZN(n5351) );
  XOR2_X2 U7302 ( .A(n5350), .B(n5349), .Z(n5375) );
  XNOR2_X2 U7303 ( .A(n5290), .B(n5289), .ZN(n5349) );
  NAND2_X2 U7305 ( .A1(n5291), .A2(n5383), .ZN(n5290) );
  OR3_X2 U7307 ( .A1(n13162), .A2(n13790), .A3(n5384), .ZN(n5291) );
  XNOR2_X2 U7308 ( .A(n5295), .B(n5294), .ZN(n5384) );
  NAND2_X2 U7310 ( .A1(n5296), .A2(n5388), .ZN(n5295) );
  OR3_X2 U7312 ( .A1(n3130), .A2(n8738), .A3(n5389), .ZN(n5296) );
  XNOR2_X2 U7313 ( .A(n5300), .B(n5299), .ZN(n5389) );
  AND3_X2 U7317 ( .A1(n13161), .A2(n13119), .A3(n5394), .ZN(n5301) );
  XOR2_X2 U7318 ( .A(n5305), .B(n5304), .Z(n5394) );
  AND3_X2 U7322 ( .A1(n13156), .A2(execstage_BusA[6]), .A3(n5399), .ZN(n5306)
         );
  XOR2_X2 U7323 ( .A(n5312), .B(n16326), .Z(n5399) );
  NAND2_X2 U7326 ( .A1(n5313), .A2(n5404), .ZN(n5312) );
  OR3_X2 U7328 ( .A1(n13215), .A2(n13155), .A3(n5405), .ZN(n5313) );
  XOR2_X2 U7329 ( .A(n5348), .B(n5346), .Z(n5405) );
  NAND2_X2 U7330 ( .A1(n5347), .A2(n5406), .ZN(n5346) );
  OR3_X2 U7332 ( .A1(n13148), .A2(n13212), .A3(n5407), .ZN(n5347) );
  XNOR2_X2 U7333 ( .A(n5341), .B(n5342), .ZN(n5407) );
  AND3_X2 U7336 ( .A1(n8648), .A2(n13211), .A3(n5409), .ZN(n5343) );
  XOR2_X2 U7337 ( .A(n5338), .B(n5339), .Z(n5409) );
  AND3_X2 U7340 ( .A1(n8694), .A2(n13207), .A3(n5411), .ZN(n5340) );
  XOR2_X2 U7341 ( .A(n5335), .B(n5336), .Z(n5411) );
  AND3_X2 U7344 ( .A1(n8652), .A2(n13188), .A3(n5413), .ZN(n5337) );
  XOR2_X2 U7345 ( .A(n5332), .B(n5333), .Z(n5413) );
  AND3_X2 U7348 ( .A1(execstage_BusA[12]), .A2(n13204), .A3(n5415), .ZN(n5334)
         );
  XOR2_X2 U7349 ( .A(n5329), .B(n5330), .Z(n5415) );
  NAND2_X2 U7355 ( .A1(n5419), .A2(n5420), .ZN(n5328) );
  XOR2_X2 U7357 ( .A(n5327), .B(n5326), .Z(n5419) );
  NAND2_X2 U7358 ( .A1(execstage_BusA[14]), .A2(n13198), .ZN(n5327) );
  NAND2_X2 U7365 ( .A1(n13166), .A2(n13792), .ZN(n5350) );
  OAI221_X2 U7369 ( .B1(n2784), .B2(n5160), .C1(n16495), .C2(n13104), .A(n5443), .ZN(n2911) );
  AOI22_X2 U7370 ( .A1(n8659), .A2(n3804), .B1(n16471), .B2(n4405), .ZN(n5443)
         );
  OAI221_X2 U7371 ( .B1(n8710), .B2(n13185), .C1(n8645), .C2(n3434), .A(n5444), 
        .ZN(n3804) );
  AOI22_X2 U7372 ( .A1(n16523), .A2(n13196), .B1(n16522), .B2(n13200), .ZN(
        n5444) );
  XOR2_X2 U7375 ( .A(n5356), .B(n5357), .Z(n5446) );
  XOR2_X2 U7376 ( .A(execstage_BusA[15]), .B(n5355), .Z(n5357) );
  XNOR2_X2 U7377 ( .A(n13133), .B(n13168), .ZN(n5355) );
  OAI22_X2 U7378 ( .A1(n16360), .A2(n8657), .B1(n5449), .B2(n5450), .ZN(n5356)
         );
  NAND4_X2 U7381 ( .A1(n5452), .A2(n5453), .A3(n5454), .A4(n5455), .ZN(
        aluout_0[14]) );
  AND3_X2 U7383 ( .A1(n5371), .A2(n13179), .A3(n8807), .ZN(n5458) );
  OAI22_X2 U7384 ( .A1(n16519), .A2(n5459), .B1(n5460), .B2(n5371), .ZN(n5456)
         );
  XNOR2_X2 U7385 ( .A(n5378), .B(n5377), .ZN(n5371) );
  NAND2_X2 U7387 ( .A1(n5379), .A2(n5462), .ZN(n5378) );
  OR3_X2 U7389 ( .A1(n13165), .A2(n13151), .A3(n5463), .ZN(n5379) );
  XNOR2_X2 U7390 ( .A(n5381), .B(n5380), .ZN(n5463) );
  AND3_X2 U7394 ( .A1(n13164), .A2(n13792), .A3(n5468), .ZN(n5382) );
  XOR2_X2 U7395 ( .A(n5385), .B(n5386), .Z(n5468) );
  AND3_X2 U7398 ( .A1(n13182), .A2(n13791), .A3(n5470), .ZN(n5387) );
  XOR2_X2 U7399 ( .A(n5391), .B(n5390), .Z(n5470) );
  NAND2_X2 U7401 ( .A1(n5392), .A2(n5474), .ZN(n5391) );
  OR3_X2 U7403 ( .A1(n13159), .A2(n8738), .A3(n5475), .ZN(n5392) );
  XNOR2_X2 U7404 ( .A(n5396), .B(n16315), .ZN(n5475) );
  NAND2_X2 U7407 ( .A1(n5397), .A2(n5480), .ZN(n5396) );
  OR3_X2 U7409 ( .A1(n13157), .A2(n13144), .A3(n5481), .ZN(n5397) );
  XNOR2_X2 U7410 ( .A(n5402), .B(n16327), .ZN(n5481) );
  NAND2_X2 U7413 ( .A1(n5403), .A2(n5486), .ZN(n5402) );
  OR3_X2 U7415 ( .A1(n13215), .A2(n13154), .A3(n5487), .ZN(n5403) );
  NAND2_X2 U7417 ( .A1(n5488), .A2(n5489), .ZN(n5441) );
  XOR2_X2 U7419 ( .A(n5439), .B(n5440), .Z(n5488) );
  XNOR2_X2 U7420 ( .A(n5436), .B(n5437), .ZN(n5439) );
  NAND2_X2 U7421 ( .A1(n5438), .A2(n5493), .ZN(n5437) );
  OR3_X2 U7423 ( .A1(n13148), .A2(n13209), .A3(n5494), .ZN(n5438) );
  XNOR2_X2 U7424 ( .A(n5433), .B(n5434), .ZN(n5494) );
  NAND2_X2 U7425 ( .A1(n5435), .A2(n5495), .ZN(n5434) );
  OR3_X2 U7427 ( .A1(n13146), .A2(n13205), .A3(n5496), .ZN(n5435) );
  XNOR2_X2 U7428 ( .A(n5430), .B(n5431), .ZN(n5496) );
  NAND2_X2 U7429 ( .A1(n5432), .A2(n5497), .ZN(n5431) );
  OR3_X2 U7431 ( .A1(n13136), .A2(n13190), .A3(n5498), .ZN(n5432) );
  XNOR2_X2 U7432 ( .A(n5427), .B(n5428), .ZN(n5498) );
  NAND2_X2 U7433 ( .A1(n5429), .A2(n5499), .ZN(n5428) );
  OR3_X2 U7435 ( .A1(n8736), .A2(n13201), .A3(n5500), .ZN(n5429) );
  XNOR2_X2 U7436 ( .A(n5424), .B(n5425), .ZN(n5500) );
  NAND2_X2 U7437 ( .A1(n5426), .A2(n5501), .ZN(n5425) );
  OR3_X2 U7439 ( .A1(n8695), .A2(n13174), .A3(n5502), .ZN(n5426) );
  NAND2_X2 U7441 ( .A1(n5503), .A2(n5504), .ZN(n5423) );
  XOR2_X2 U7443 ( .A(n5422), .B(n5421), .Z(n5503) );
  NAND2_X2 U7444 ( .A1(n13120), .A2(n13199), .ZN(n5422) );
  AOI221_X2 U7454 ( .B1(n2726), .B2(n4667), .C1(n16456), .C2(n3234), .A(n16399), .ZN(n5453) );
  AOI22_X2 U7456 ( .A1(n4668), .A2(n2724), .B1(n2805), .B2(n16449), .ZN(n5528)
         );
  OAI221_X2 U7457 ( .B1(n16513), .B2(n5160), .C1(n16514), .C2(n13104), .A(
        n5529), .ZN(n3234) );
  AOI22_X2 U7458 ( .A1(n8659), .A2(n3965), .B1(n16471), .B2(n5071), .ZN(n5529)
         );
  OAI221_X2 U7459 ( .B1(n13137), .B2(n13184), .C1(n8657), .C2(n3434), .A(n5530), .ZN(n3965) );
  AOI22_X2 U7460 ( .A1(n16542), .A2(n13200), .B1(n16543), .B2(n13195), .ZN(
        n5530) );
  XOR2_X2 U7463 ( .A(n5450), .B(n5449), .Z(n5533) );
  AOI22_X2 U7464 ( .A1(n5536), .A2(n8655), .B1(n5537), .B2(n5538), .ZN(n5449)
         );
  XOR2_X2 U7465 ( .A(n13138), .B(n5451), .Z(n5450) );
  XNOR2_X2 U7466 ( .A(n13133), .B(n13179), .ZN(n5451) );
  NAND4_X2 U7468 ( .A1(n5539), .A2(n5540), .A3(n5541), .A4(n5542), .ZN(
        aluout_0[13]) );
  OAI22_X2 U7472 ( .A1(n16517), .A2(n5459), .B1(n5546), .B2(n5545), .ZN(n5543)
         );
  XNOR2_X2 U7473 ( .A(n5465), .B(n5464), .ZN(n5545) );
  NAND2_X2 U7475 ( .A1(n5466), .A2(n5548), .ZN(n5465) );
  OR3_X2 U7477 ( .A1(n13162), .A2(n13151), .A3(n5549), .ZN(n5466) );
  NAND2_X2 U7479 ( .A1(n5550), .A2(n5551), .ZN(n5525) );
  XOR2_X2 U7481 ( .A(n5524), .B(n5523), .Z(n5550) );
  XNOR2_X2 U7482 ( .A(n5472), .B(n5471), .ZN(n5523) );
  AND3_X2 U7486 ( .A1(n13161), .A2(n13791), .A3(n5559), .ZN(n5473) );
  XOR2_X2 U7487 ( .A(n5478), .B(n5477), .Z(n5559) );
  NAND2_X2 U7489 ( .A1(n5479), .A2(n5563), .ZN(n5478) );
  OR3_X2 U7491 ( .A1(n13157), .A2(n8738), .A3(n5564), .ZN(n5479) );
  XNOR2_X2 U7492 ( .A(n5484), .B(n16328), .ZN(n5564) );
  NAND2_X2 U7495 ( .A1(n5485), .A2(n5569), .ZN(n5484) );
  OR3_X2 U7497 ( .A1(n13215), .A2(n13144), .A3(n5570), .ZN(n5485) );
  XNOR2_X2 U7498 ( .A(n5491), .B(n16340), .ZN(n5570) );
  NAND2_X2 U7501 ( .A1(n5492), .A2(n5575), .ZN(n5491) );
  OR3_X2 U7503 ( .A1(n13212), .A2(n8715), .A3(n5576), .ZN(n5492) );
  XNOR2_X2 U7504 ( .A(n5520), .B(n5521), .ZN(n5576) );
  AND3_X2 U7507 ( .A1(execstage_BusA[7]), .A2(n13211), .A3(n5578), .ZN(n5522)
         );
  XOR2_X2 U7508 ( .A(n5517), .B(n5518), .Z(n5578) );
  AND3_X2 U7511 ( .A1(execstage_BusA[8]), .A2(n13207), .A3(n5580), .ZN(n5519)
         );
  XOR2_X2 U7512 ( .A(n5514), .B(n5515), .Z(n5580) );
  AND3_X2 U7515 ( .A1(n8648), .A2(n13188), .A3(n5582), .ZN(n5516) );
  XOR2_X2 U7516 ( .A(n5511), .B(n5512), .Z(n5582) );
  AND3_X2 U7519 ( .A1(n8694), .A2(n13204), .A3(n5584), .ZN(n5513) );
  XOR2_X2 U7520 ( .A(n5508), .B(n5509), .Z(n5584) );
  NAND2_X2 U7526 ( .A1(n5588), .A2(n5589), .ZN(n5507) );
  XOR2_X2 U7528 ( .A(n5506), .B(n5505), .Z(n5588) );
  NAND2_X2 U7529 ( .A1(execstage_BusA[12]), .A2(n13198), .ZN(n5506) );
  NAND2_X2 U7535 ( .A1(n13182), .A2(n13792), .ZN(n5524) );
  AOI22_X2 U7542 ( .A1(n13171), .A2(execstage_BusA[29]), .B1(n13194), .B2(
        n2921), .ZN(n5608) );
  AOI22_X2 U7545 ( .A1(n5240), .A2(n5264), .B1(n16523), .B2(n13195), .ZN(n5612) );
  NAND2_X2 U7547 ( .A1(n5239), .A2(n13198), .ZN(n5054) );
  AOI221_X2 U7548 ( .B1(n2726), .B2(n4246), .C1(n16456), .C2(n3430), .A(n16396), .ZN(n5540) );
  AOI22_X2 U7550 ( .A1(n2727), .A2(n2724), .B1(n2725), .B2(n16449), .ZN(n5614)
         );
  OAI211_X2 U7551 ( .C1(n13194), .C2(n4766), .A(n5261), .B(n5615), .ZN(n2725)
         );
  AOI22_X2 U7552 ( .A1(n5616), .A2(n13196), .B1(execstage_BusA[19]), .B2(
        n13183), .ZN(n5615) );
  NAND2_X2 U7553 ( .A1(execstage_BusA[17]), .A2(n13171), .ZN(n5261) );
  OAI221_X2 U7554 ( .B1(n13185), .B2(n8656), .C1(n13169), .C2(n8646), .A(n5617), .ZN(n2727) );
  AOI22_X2 U7555 ( .A1(n16526), .A2(n13196), .B1(n16527), .B2(n13200), .ZN(
        n5617) );
  OAI221_X2 U7556 ( .B1(n16491), .B2(n13103), .C1(n16490), .C2(n2873), .A(
        n5618), .ZN(n3430) );
  AOI22_X2 U7557 ( .A1(n8696), .A2(n2839), .B1(n16469), .B2(n4941), .ZN(n5618)
         );
  NAND2_X2 U7559 ( .A1(n13171), .A2(execstage_BusA[1]), .ZN(n4933) );
  OAI221_X2 U7560 ( .B1(n13790), .B2(n13184), .C1(n13143), .C2(n3434), .A(
        n5620), .ZN(n2839) );
  AOI22_X2 U7561 ( .A1(n16530), .A2(n13196), .B1(n4931), .B2(n13197), .ZN(
        n5620) );
  OAI221_X2 U7563 ( .B1(n13155), .B2(n13184), .C1(n13146), .C2(n3434), .A(
        n5622), .ZN(n5174) );
  AOI22_X2 U7564 ( .A1(n16532), .A2(n13196), .B1(n16531), .B2(n13197), .ZN(
        n5622) );
  OAI211_X2 U7566 ( .C1(n13197), .C2(n5590), .A(n5611), .B(n5625), .ZN(n4683)
         );
  AOI22_X2 U7567 ( .A1(n16529), .A2(n13198), .B1(n13183), .B2(n8652), .ZN(
        n5625) );
  NAND2_X2 U7568 ( .A1(n13171), .A2(n8655), .ZN(n5611) );
  OAI221_X2 U7569 ( .B1(n13185), .B2(n8713), .C1(n13169), .C2(n8732), .A(n5626), .ZN(n4246) );
  AOI22_X2 U7570 ( .A1(n16528), .A2(n13196), .B1(n16524), .B2(n13200), .ZN(
        n5626) );
  XOR2_X2 U7572 ( .A(n5537), .B(n5538), .Z(n5628) );
  XOR2_X2 U7573 ( .A(n8655), .B(n5536), .Z(n5538) );
  XNOR2_X2 U7574 ( .A(n13133), .B(n13166), .ZN(n5536) );
  OAI22_X2 U7575 ( .A1(n16365), .A2(n8695), .B1(n5631), .B2(n5632), .ZN(n5537)
         );
  NAND4_X2 U7578 ( .A1(n5634), .A2(n5635), .A3(n5636), .A4(n5637), .ZN(
        aluout_0[12]) );
  AOI22_X2 U7584 ( .A1(n4387), .A2(n13174), .B1(n13177), .B2(n4388), .ZN(n2851) );
  AOI22_X2 U7586 ( .A1(n4928), .A2(n13198), .B1(n16545), .B2(n13195), .ZN(
        n5645) );
  AOI221_X2 U7588 ( .B1(n5547), .B2(n5647), .C1(n13218), .C2(n5648), .A(n16402), .ZN(n5636) );
  AOI22_X2 U7590 ( .A1(n2749), .A2(n16449), .B1(n2751), .B2(n16448), .ZN(n5650) );
  XOR2_X2 U7592 ( .A(n5553), .B(n5552), .Z(n5547) );
  NAND2_X2 U7594 ( .A1(n5554), .A2(n5652), .ZN(n5553) );
  OR3_X2 U7596 ( .A1(n3130), .A2(n13151), .A3(n5653), .ZN(n5554) );
  XNOR2_X2 U7597 ( .A(n5556), .B(n5555), .ZN(n5653) );
  NAND2_X2 U7599 ( .A1(n5557), .A2(n5657), .ZN(n5556) );
  OR3_X2 U7601 ( .A1(n13159), .A2(n13793), .A3(n5658), .ZN(n5557) );
  XNOR2_X2 U7602 ( .A(n5560), .B(n5561), .ZN(n5658) );
  AND3_X2 U7605 ( .A1(n13156), .A2(n13791), .A3(n5660), .ZN(n5562) );
  XOR2_X2 U7606 ( .A(n5567), .B(n5566), .Z(n5660) );
  NAND2_X2 U7608 ( .A1(n5568), .A2(n5664), .ZN(n5567) );
  OR3_X2 U7610 ( .A1(n13215), .A2(n8738), .A3(n5665), .ZN(n5568) );
  XNOR2_X2 U7611 ( .A(n5573), .B(n16341), .ZN(n5665) );
  NAND2_X2 U7614 ( .A1(n5574), .A2(n5670), .ZN(n5573) );
  OR3_X2 U7616 ( .A1(n13212), .A2(n13144), .A3(n5671), .ZN(n5574) );
  NAND2_X2 U7618 ( .A1(n5672), .A2(n5673), .ZN(n5607) );
  XOR2_X2 U7620 ( .A(n5605), .B(n5606), .Z(n5672) );
  XNOR2_X2 U7621 ( .A(n5602), .B(n5603), .ZN(n5605) );
  NAND2_X2 U7622 ( .A1(n5604), .A2(n5677), .ZN(n5603) );
  OR3_X2 U7624 ( .A1(n13155), .A2(n13205), .A3(n5678), .ZN(n5604) );
  XNOR2_X2 U7625 ( .A(n5599), .B(n5600), .ZN(n5678) );
  NAND2_X2 U7626 ( .A1(n5601), .A2(n5679), .ZN(n5600) );
  OR3_X2 U7628 ( .A1(n13148), .A2(n13190), .A3(n5680), .ZN(n5601) );
  XNOR2_X2 U7629 ( .A(n5596), .B(n5597), .ZN(n5680) );
  NAND2_X2 U7630 ( .A1(n5598), .A2(n5681), .ZN(n5597) );
  OR3_X2 U7632 ( .A1(n13146), .A2(n13201), .A3(n5682), .ZN(n5598) );
  XNOR2_X2 U7633 ( .A(n5594), .B(n16475), .ZN(n5682) );
  NAND2_X2 U7637 ( .A1(n5595), .A2(n5688), .ZN(n5594) );
  OR3_X2 U7639 ( .A1(n13136), .A2(n13174), .A3(n5689), .ZN(n5595) );
  NAND2_X2 U7641 ( .A1(n5690), .A2(n5691), .ZN(n5592) );
  XOR2_X2 U7643 ( .A(n5591), .B(n5590), .Z(n5690) );
  NAND2_X2 U7644 ( .A1(n13121), .A2(n13199), .ZN(n5591) );
  AOI221_X2 U7649 ( .B1(n2724), .B2(n2753), .C1(n2726), .C2(n4261), .A(n16454), 
        .ZN(n5635) );
  AOI22_X2 U7651 ( .A1(n3643), .A2(n13106), .B1(n3645), .B2(n16455), .ZN(n5708) );
  OAI221_X2 U7652 ( .B1(n13154), .B2(n13184), .C1(n13148), .C2(n13169), .A(
        n5709), .ZN(n3645) );
  AOI22_X2 U7653 ( .A1(n16540), .A2(n13196), .B1(n16539), .B2(n13200), .ZN(
        n5709) );
  OAI221_X2 U7654 ( .B1(n13136), .B2(n13184), .C1(n13137), .C2(n13170), .A(
        n5712), .ZN(n3643) );
  AOI22_X2 U7655 ( .A1(n16542), .A2(n13196), .B1(n16541), .B2(n13200), .ZN(
        n5712) );
  XOR2_X2 U7658 ( .A(n5632), .B(n5631), .Z(n5715) );
  AOI22_X2 U7659 ( .A1(n5718), .A2(n8652), .B1(n5719), .B2(n5720), .ZN(n5631)
         );
  XOR2_X2 U7660 ( .A(n13137), .B(n5633), .Z(n5632) );
  XNOR2_X2 U7661 ( .A(n13134), .B(n13164), .ZN(n5633) );
  NAND4_X2 U7663 ( .A1(n5721), .A2(n5722), .A3(n16370), .A4(n5724), .ZN(
        aluout_0[11]) );
  AOI221_X2 U7664 ( .B1(n5725), .B2(n5726), .C1(n16317), .C2(n5727), .A(n5728), 
        .ZN(n5724) );
  NAND2_X2 U7666 ( .A1(n16458), .A2(n13103), .ZN(n5641) );
  NAND2_X2 U7668 ( .A1(execstage_ALU_ra_row2_31_), .A2(n2733), .ZN(n3954) );
  NAND2_X2 U7669 ( .A1(n13114), .A2(n13201), .ZN(n5729) );
  OAI22_X2 U7670 ( .A1(n13177), .A2(n3803), .B1(n16518), .B2(n13174), .ZN(
        n3801) );
  NAND2_X2 U7672 ( .A1(n13171), .A2(execstage_ALU_ra_row2_31_), .ZN(n4530) );
  XNOR2_X2 U7675 ( .A(n5655), .B(n5654), .ZN(n5726) );
  NAND2_X2 U7682 ( .A1(n5734), .A2(n5735), .ZN(n5706) );
  XOR2_X2 U7684 ( .A(n5705), .B(n5704), .Z(n5734) );
  XNOR2_X2 U7685 ( .A(n5662), .B(n5661), .ZN(n5704) );
  AND3_X2 U7689 ( .A1(n13217), .A2(n13791), .A3(n5743), .ZN(n5663) );
  XOR2_X2 U7690 ( .A(n5668), .B(n16342), .Z(n5743) );
  NAND2_X2 U7693 ( .A1(n5669), .A2(n5748), .ZN(n5668) );
  OR3_X2 U7695 ( .A1(n13212), .A2(n8738), .A3(n5749), .ZN(n5669) );
  XNOR2_X2 U7696 ( .A(n5675), .B(n16343), .ZN(n5749) );
  NAND2_X2 U7699 ( .A1(n5676), .A2(n5754), .ZN(n5675) );
  OR3_X2 U7701 ( .A1(n13209), .A2(n13143), .A3(n5755), .ZN(n5676) );
  XNOR2_X2 U7702 ( .A(n5701), .B(n5702), .ZN(n5755) );
  AND3_X2 U7705 ( .A1(execstage_BusA[6]), .A2(n13208), .A3(n5757), .ZN(n5703)
         );
  XOR2_X2 U7706 ( .A(n5698), .B(n5699), .Z(n5757) );
  AND3_X2 U7709 ( .A1(n13115), .A2(n13188), .A3(n5759), .ZN(n5700) );
  XOR2_X2 U7710 ( .A(n5695), .B(n5696), .Z(n5759) );
  AND3_X2 U7713 ( .A1(execstage_BusA[8]), .A2(n13204), .A3(n5761), .ZN(n5697)
         );
  XNOR2_X2 U7714 ( .A(n5687), .B(n5685), .ZN(n5761) );
  NAND2_X2 U7715 ( .A1(n5686), .A2(n5762), .ZN(n5685) );
  OR3_X2 U7717 ( .A1(n13146), .A2(n13175), .A3(n5763), .ZN(n5686) );
  NAND2_X2 U7719 ( .A1(n5764), .A2(n5765), .ZN(n5694) );
  XOR2_X2 U7721 ( .A(n5693), .B(n5692), .Z(n5764) );
  NAND2_X2 U7722 ( .A1(n13122), .A2(n13199), .ZN(n5693) );
  NAND2_X2 U7727 ( .A1(n13158), .A2(n13792), .ZN(n5705) );
  OAI221_X2 U7730 ( .B1(n5459), .B2(n16494), .C1(n13220), .C2(n5781), .A(n5782), .ZN(n5780) );
  AOI22_X2 U7731 ( .A1(n2777), .A2(n16448), .B1(n16509), .B2(n3807), .ZN(n5782) );
  AOI221_X2 U7734 ( .B1(n13194), .B2(n4931), .C1(execstage_BusA[1]), .C2(
        n13183), .A(n5783), .ZN(n2784) );
  OAI22_X2 U7735 ( .A1(n13170), .A2(n13790), .B1(n5619), .B2(n13196), .ZN(
        n5783) );
  OAI221_X2 U7736 ( .B1(n8710), .B2(n13184), .C1(n8736), .C2(n13169), .A(n5784), .ZN(n2777) );
  AOI22_X2 U7737 ( .A1(n16523), .A2(n13198), .B1(n16522), .B2(n13195), .ZN(
        n5784) );
  NAND2_X2 U7739 ( .A1(execstage_BusA[12]), .A2(n13129), .ZN(n5590) );
  NAND2_X2 U7741 ( .A1(execstage_BusA[14]), .A2(n13129), .ZN(n5421) );
  OAI221_X2 U7743 ( .B1(n13185), .B2(n8737), .C1(n13169), .C2(n8713), .A(n5785), .ZN(n3803) );
  AOI22_X2 U7744 ( .A1(n2921), .A2(n13198), .B1(n16524), .B2(n13195), .ZN(
        n5785) );
  NAND2_X2 U7746 ( .A1(execstage_BusA[28]), .A2(n13129), .ZN(n2917) );
  NAND2_X2 U7748 ( .A1(n8659), .A2(n2733), .ZN(n5459) );
  AOI221_X2 U7749 ( .B1(n2726), .B2(n4531), .C1(n16455), .C2(n2790), .A(n16386), .ZN(n5722) );
  AOI22_X2 U7751 ( .A1(n2776), .A2(n2724), .B1(n2778), .B2(n16449), .ZN(n5787)
         );
  OAI221_X2 U7752 ( .B1(n13185), .B2(n8647), .C1(n8645), .C2(n13169), .A(n5788), .ZN(n2778) );
  NAND2_X2 U7758 ( .A1(n5239), .A2(n13196), .ZN(n5262) );
  OAI221_X2 U7760 ( .B1(n13185), .B2(n8646), .C1(n13169), .C2(n8654), .A(n5790), .ZN(n2776) );
  AOI22_X2 U7761 ( .A1(n16526), .A2(n13198), .B1(n16525), .B2(n13195), .ZN(
        n5790) );
  NAND2_X2 U7763 ( .A1(execstage_BusA[20]), .A2(n13129), .ZN(n4766) );
  NAND2_X2 U7765 ( .A1(execstage_BusA[22]), .A2(n13129), .ZN(n4492) );
  OAI221_X2 U7766 ( .B1(n13143), .B2(n13184), .C1(n13155), .C2(n13169), .A(
        n5791), .ZN(n2790) );
  AOI22_X2 U7767 ( .A1(n16531), .A2(n13196), .B1(n16530), .B2(n13200), .ZN(
        n5791) );
  NAND2_X2 U7771 ( .A1(n16471), .A2(n16456), .ZN(n2785) );
  OAI221_X2 U7772 ( .B1(n13185), .B2(n8732), .C1(n13169), .C2(n8656), .A(n5792), .ZN(n4531) );
  AOI22_X2 U7773 ( .A1(n16528), .A2(n13198), .B1(n16527), .B2(n13195), .ZN(
        n5792) );
  NAND2_X2 U7775 ( .A1(execstage_BusA[24]), .A2(n13129), .ZN(n4206) );
  NAND2_X2 U7777 ( .A1(execstage_BusA[26]), .A2(n13129), .ZN(n3908) );
  AOI221_X2 U7778 ( .B1(n13106), .B2(n4405), .C1(n5793), .C2(n13783), .A(
        n16368), .ZN(n5721) );
  AOI22_X2 U7780 ( .A1(n16548), .A2(n16369), .B1(n13130), .B2(n5796), .ZN(
        n5795) );
  XOR2_X2 U7781 ( .A(n5719), .B(n5720), .Z(n5793) );
  XOR2_X2 U7782 ( .A(n8652), .B(n5718), .Z(n5720) );
  XNOR2_X2 U7783 ( .A(n13134), .B(n13182), .ZN(n5718) );
  OAI22_X2 U7784 ( .A1(n16416), .A2(n13136), .B1(n5798), .B2(n5799), .ZN(n5719) );
  OAI221_X2 U7786 ( .B1(n13146), .B2(n13184), .C1(n8736), .C2(n13169), .A(
        n5801), .ZN(n4405) );
  AOI22_X2 U7787 ( .A1(n16529), .A2(n13195), .B1(n16532), .B2(n13200), .ZN(
        n5801) );
  NAND4_X2 U7790 ( .A1(n5802), .A2(n5803), .A3(n5804), .A4(n5805), .ZN(
        aluout_0[10]) );
  AOI221_X2 U7791 ( .B1(n5806), .B2(n5730), .C1(n16320), .C2(n5808), .A(n5809), 
        .ZN(n5805) );
  OAI22_X2 U7792 ( .A1(n5810), .A2(n13220), .B1(n3962), .B2(n8722), .ZN(n5809)
         );
  AOI22_X2 U7795 ( .A1(n4667), .A2(n8659), .B1(n3247), .B2(n16471), .ZN(n3962)
         );
  NAND2_X2 U7796 ( .A1(n5811), .A2(n3243), .ZN(n3247) );
  NAND2_X2 U7799 ( .A1(n8649), .A2(n8712), .ZN(n2715) );
  XNOR2_X2 U7801 ( .A(n5737), .B(n5736), .ZN(n5730) );
  XOR2_X2 U7803 ( .A(n5812), .B(n5813), .Z(n2707) );
  NAND2_X2 U7804 ( .A1(n5738), .A2(n5814), .ZN(n5737) );
  OR3_X2 U7806 ( .A1(n13157), .A2(n13151), .A3(n5815), .ZN(n5738) );
  XNOR2_X2 U7807 ( .A(n5740), .B(n5739), .ZN(n5815) );
  XNOR2_X2 U7815 ( .A(n5823), .B(n5824), .ZN(n2740) );
  NAND2_X2 U7816 ( .A1(n5741), .A2(n5825), .ZN(n5740) );
  OR3_X2 U7818 ( .A1(n13215), .A2(n13793), .A3(n5826), .ZN(n5741) );
  XNOR2_X2 U7819 ( .A(n5746), .B(n16345), .ZN(n5826) );
  NAND2_X2 U7822 ( .A1(n5820), .A2(n5821), .ZN(n5822) );
  NAND2_X2 U7824 ( .A1(n5830), .A2(n5831), .ZN(n5823) );
  OR3_X2 U7826 ( .A1(n13212), .A2(n13151), .A3(n5832), .ZN(n5830) );
  XNOR2_X2 U7827 ( .A(n5833), .B(n5834), .ZN(n5832) );
  XNOR2_X2 U7830 ( .A(n5835), .B(n5836), .ZN(n2767) );
  XOR2_X2 U7831 ( .A(n5829), .B(n5828), .Z(n5820) );
  NAND2_X2 U7832 ( .A1(n13214), .A2(n13792), .ZN(n5829) );
  XNOR2_X2 U7833 ( .A(n5837), .B(n5838), .ZN(n5828) );
  NAND2_X2 U7834 ( .A1(n5747), .A2(n5839), .ZN(n5746) );
  OR3_X2 U7836 ( .A1(n13212), .A2(n13790), .A3(n5840), .ZN(n5747) );
  XNOR2_X2 U7837 ( .A(n5752), .B(n5751), .ZN(n5840) );
  XOR2_X2 U7843 ( .A(n5845), .B(n5846), .Z(n5844) );
  NAND2_X2 U7845 ( .A1(n5847), .A2(n5848), .ZN(n5833) );
  OR3_X2 U7847 ( .A1(n13209), .A2(n13793), .A3(n5849), .ZN(n5847) );
  XNOR2_X2 U7848 ( .A(n5850), .B(n5851), .ZN(n5849) );
  XNOR2_X2 U7856 ( .A(n5859), .B(n5860), .ZN(n2797) );
  NAND2_X2 U7857 ( .A1(n5753), .A2(n5861), .ZN(n5752) );
  OR3_X2 U7859 ( .A1(n13209), .A2(n8738), .A3(n5862), .ZN(n5753) );
  NAND2_X2 U7861 ( .A1(n5863), .A2(n5864), .ZN(n5779) );
  NAND2_X2 U7863 ( .A1(n5866), .A2(n5867), .ZN(n5846) );
  OR3_X2 U7865 ( .A1(n13205), .A2(n8738), .A3(n5868), .ZN(n5866) );
  XNOR2_X2 U7866 ( .A(n5869), .B(n5870), .ZN(n5868) );
  NAND2_X2 U7869 ( .A1(n5871), .A2(n5872), .ZN(n5850) );
  OR3_X2 U7871 ( .A1(n13205), .A2(n13790), .A3(n5873), .ZN(n5871) );
  NAND2_X2 U7875 ( .A1(n5856), .A2(n5857), .ZN(n5858) );
  NAND2_X2 U7877 ( .A1(n5880), .A2(n5881), .ZN(n5860) );
  OR3_X2 U7879 ( .A1(n13205), .A2(n13152), .A3(n5882), .ZN(n5880) );
  XNOR2_X2 U7880 ( .A(n5883), .B(n5884), .ZN(n5882) );
  XNOR2_X2 U7883 ( .A(n5885), .B(n5886), .ZN(n2823) );
  XOR2_X2 U7884 ( .A(n5877), .B(n5878), .Z(n5856) );
  XOR2_X2 U7886 ( .A(n5887), .B(n5888), .Z(n5877) );
  XOR2_X2 U7887 ( .A(n5777), .B(n5778), .Z(n5863) );
  XNOR2_X2 U7888 ( .A(n5774), .B(n5775), .ZN(n5777) );
  NAND2_X2 U7889 ( .A1(n5776), .A2(n5889), .ZN(n5775) );
  OR3_X2 U7891 ( .A1(n13154), .A2(n13190), .A3(n5890), .ZN(n5776) );
  XNOR2_X2 U7892 ( .A(n5771), .B(n5772), .ZN(n5890) );
  NAND2_X2 U7893 ( .A1(n5773), .A2(n5891), .ZN(n5772) );
  OR3_X2 U7895 ( .A1(n13155), .A2(n13201), .A3(n5892), .ZN(n5773) );
  XNOR2_X2 U7896 ( .A(n5769), .B(n16477), .ZN(n5892) );
  NAND2_X2 U7904 ( .A1(n5900), .A2(n5901), .ZN(n5767) );
  XOR2_X2 U7906 ( .A(n5766), .B(n2884), .Z(n5900) );
  NAND2_X2 U7907 ( .A1(n8694), .A2(n13129), .ZN(n2884) );
  NAND2_X2 U7908 ( .A1(n13118), .A2(n13199), .ZN(n5766) );
  AND3_X2 U7913 ( .A1(n13119), .A2(n13188), .A3(n5909), .ZN(n5907) );
  XOR2_X2 U7914 ( .A(n5904), .B(n5905), .Z(n5909) );
  AND3_X2 U7917 ( .A1(n13116), .A2(n13204), .A3(n5911), .ZN(n5906) );
  XOR2_X2 U7918 ( .A(n5895), .B(n5894), .Z(n5911) );
  NAND2_X2 U7925 ( .A1(n5918), .A2(n5919), .ZN(n5903) );
  XOR2_X2 U7927 ( .A(n5902), .B(n3411), .Z(n5918) );
  NAND2_X2 U7928 ( .A1(execstage_BusA[8]), .A2(n13199), .ZN(n5902) );
  NAND2_X2 U7931 ( .A1(n5874), .A2(n5875), .ZN(n5876) );
  NAND2_X2 U7933 ( .A1(n5926), .A2(n5927), .ZN(n5888) );
  OR3_X2 U7935 ( .A1(n13790), .A2(n13190), .A3(n5928), .ZN(n5926) );
  XNOR2_X2 U7936 ( .A(n5929), .B(n5930), .ZN(n5928) );
  NAND2_X2 U7944 ( .A1(n5938), .A2(n5939), .ZN(n5885) );
  OR3_X2 U7946 ( .A1(n13151), .A2(n13190), .A3(n5940), .ZN(n5938) );
  XOR2_X2 U7949 ( .A(n5944), .B(n5945), .Z(n2845) );
  XOR2_X2 U7950 ( .A(n2861), .B(n5925), .Z(n5874) );
  XNOR2_X2 U7951 ( .A(n5923), .B(n5922), .ZN(n5925) );
  AND3_X2 U7955 ( .A1(execstage_BusA[4]), .A2(n13204), .A3(n5948), .ZN(n5946)
         );
  XOR2_X2 U7956 ( .A(n5949), .B(n5950), .Z(n5948) );
  NAND2_X2 U7958 ( .A1(n5935), .A2(n5936), .ZN(n5937) );
  NAND2_X2 U7960 ( .A1(n5941), .A2(n5942), .ZN(n5943) );
  NAND2_X2 U7962 ( .A1(n5954), .A2(n5955), .ZN(n5945) );
  OR3_X2 U7964 ( .A1(n13201), .A2(n13152), .A3(n5956), .ZN(n5954) );
  XNOR2_X2 U7965 ( .A(n5957), .B(n5958), .ZN(n5956) );
  XOR2_X2 U7967 ( .A(n5959), .B(n5960), .Z(n2866) );
  XOR2_X2 U7968 ( .A(n5952), .B(n5953), .Z(n5941) );
  NAND2_X2 U7969 ( .A1(n13204), .A2(execstage_BusA[2]), .ZN(n5953) );
  XNOR2_X2 U7970 ( .A(n5961), .B(n5962), .ZN(n5952) );
  XOR2_X2 U7971 ( .A(n2897), .B(n5951), .Z(n5935) );
  XNOR2_X2 U7972 ( .A(n5963), .B(n5964), .ZN(n5951) );
  NAND2_X2 U7973 ( .A1(n5924), .A2(n5965), .ZN(n5923) );
  OR3_X2 U7975 ( .A1(n13143), .A2(n13201), .A3(n5966), .ZN(n5924) );
  XNOR2_X2 U7976 ( .A(n5913), .B(n5912), .ZN(n5966) );
  NAND2_X2 U7986 ( .A1(n13177), .A2(execstage_BusA[4]), .ZN(n5976) );
  AOI22_X2 U7994 ( .A1(n3421), .A2(n16501), .B1(n5957), .B2(n5958), .ZN(n5962)
         );
  XOR2_X2 U7995 ( .A(n3421), .B(n16501), .Z(n5958) );
  XOR2_X2 U7999 ( .A(n5991), .B(n5992), .Z(n5990) );
  OR3_X2 U8001 ( .A1(n8712), .A2(n3398), .A3(n13174), .ZN(n5960) );
  XNOR2_X2 U8002 ( .A(n5993), .B(n5994), .ZN(n3398) );
  XOR2_X2 U8003 ( .A(n16504), .B(n4931), .Z(n5994) );
  NAND2_X2 U8008 ( .A1(n13177), .A2(n13116), .ZN(n6000) );
  NAND2_X2 U8010 ( .A1(n6001), .A2(n6002), .ZN(n5921) );
  NAND2_X2 U8012 ( .A1(n5971), .A2(n5972), .ZN(n5973) );
  NAND2_X2 U8014 ( .A1(n5977), .A2(n5978), .ZN(n5979) );
  NAND2_X2 U8016 ( .A1(n5984), .A2(n5985), .ZN(n5986) );
  NAND2_X2 U8018 ( .A1(n5996), .A2(n5997), .ZN(n5998) );
  NAND2_X2 U8020 ( .A1(n6007), .A2(n6008), .ZN(n5992) );
  NAND2_X2 U8022 ( .A1(n6009), .A2(n13792), .ZN(n6007) );
  AND3_X2 U8024 ( .A1(n4928), .A2(n13199), .A3(execstage_BusA[0]), .ZN(n5993)
         );
  XOR2_X2 U8027 ( .A(n6006), .B(n2880), .Z(n5996) );
  NAND2_X2 U8028 ( .A1(n13791), .A2(n13199), .ZN(n6006) );
  NAND2_X2 U8029 ( .A1(execstage_BusA[4]), .A2(n13129), .ZN(n2880) );
  XOR2_X2 U8030 ( .A(n6005), .B(n3408), .Z(n5984) );
  NAND2_X2 U8031 ( .A1(execstage_BusA[4]), .A2(n13199), .ZN(n6005) );
  XOR2_X2 U8032 ( .A(n6004), .B(n2882), .Z(n5977) );
  NAND2_X2 U8033 ( .A1(n13119), .A2(n13199), .ZN(n6004) );
  NAND2_X2 U8034 ( .A1(n13116), .A2(n13129), .ZN(n2882) );
  XOR2_X2 U8035 ( .A(n6003), .B(n3412), .Z(n5971) );
  NAND2_X2 U8036 ( .A1(execstage_BusA[6]), .A2(n13199), .ZN(n6003) );
  XOR2_X2 U8037 ( .A(n5920), .B(n2885), .Z(n6001) );
  NAND2_X2 U8038 ( .A1(execstage_BusA[8]), .A2(n13129), .ZN(n2885) );
  NAND2_X2 U8039 ( .A1(execstage_BusA[7]), .A2(n13199), .ZN(n5920) );
  OAI221_X2 U8042 ( .B1(n13139), .B2(n13184), .C1(n13138), .C2(n3434), .A(
        n6011), .ZN(n2807) );
  AOI22_X2 U8043 ( .A1(n16544), .A2(n13195), .B1(n16536), .B2(n13197), .ZN(
        n6011) );
  NAND2_X2 U8045 ( .A1(n5358), .A2(n16471), .ZN(n4929) );
  OAI221_X2 U8046 ( .B1(n13137), .B2(n13184), .C1(n13136), .C2(n3434), .A(
        n6012), .ZN(n2806) );
  AOI22_X2 U8047 ( .A1(n16542), .A2(n13195), .B1(n16543), .B2(n13197), .ZN(
        n6012) );
  NAND2_X2 U8049 ( .A1(n5358), .A2(n8659), .ZN(n2772) );
  OAI221_X2 U8050 ( .B1(n13185), .B2(n13117), .C1(n13169), .C2(n8650), .A(
        n6013), .ZN(n2805) );
  NAND2_X2 U8053 ( .A1(n16535), .A2(n13199), .ZN(n4390) );
  AOI221_X2 U8057 ( .B1(n3245), .B2(n16471), .C1(n4667), .C2(n8659), .A(n16462), .ZN(n6014) );
  NAND2_X2 U8059 ( .A1(n13204), .A2(execstage_ALU_ra_row2_31_), .ZN(n4245) );
  AOI22_X2 U8061 ( .A1(n16537), .A2(n13195), .B1(n3238), .B2(n13197), .ZN(
        n6015) );
  NAND2_X2 U8062 ( .A1(execstage_BusA[28]), .A2(n13183), .ZN(n3241) );
  NAND2_X2 U8063 ( .A1(execstage_BusA[26]), .A2(n13171), .ZN(n4100) );
  NAND2_X2 U8065 ( .A1(execstage_BusA[30]), .A2(n13171), .ZN(n3243) );
  OAI221_X2 U8067 ( .B1(n13186), .B2(n8731), .C1(n13169), .C2(n8653), .A(n6017), .ZN(n4668) );
  OAI222_X2 U8073 ( .A1(n16513), .A2(n13104), .B1(n16503), .B2(n13103), .C1(
        n16514), .C2(n2873), .ZN(n4104) );
  OAI221_X2 U8075 ( .B1(n8738), .B2(n13184), .C1(n13154), .C2(n13170), .A(
        n6018), .ZN(n2816) );
  OAI221_X2 U8078 ( .B1(n13148), .B2(n13184), .C1(n13136), .C2(n13170), .A(
        n6019), .ZN(n5071) );
  AOI22_X2 U8079 ( .A1(n16541), .A2(n13195), .B1(n16540), .B2(n13197), .ZN(
        n6019) );
  OAI211_X2 U8082 ( .C1(n8712), .C2(n13185), .A(n3409), .B(n6020), .ZN(n3420)
         );
  NAND2_X2 U8083 ( .A1(n13171), .A2(execstage_BusA[2]), .ZN(n3409) );
  XOR2_X2 U8087 ( .A(n5799), .B(n5798), .Z(n6022) );
  AOI22_X2 U8088 ( .A1(n6024), .A2(n8648), .B1(n16331), .B2(n2729), .ZN(n5798)
         );
  XOR2_X2 U8089 ( .A(n13118), .B(n6024), .Z(n2729) );
  AOI22_X2 U8091 ( .A1(n6026), .A2(execstage_BusA[8]), .B1(n2756), .B2(n2755), 
        .ZN(n6025) );
  XOR2_X2 U8092 ( .A(execstage_BusA[8]), .B(n6026), .Z(n2755) );
  OAI22_X2 U8093 ( .A1(n6027), .A2(n13155), .B1(n2786), .B2(n2787), .ZN(n2756)
         );
  XOR2_X2 U8094 ( .A(n13115), .B(n6027), .Z(n2787) );
  AOI22_X2 U8095 ( .A1(n6028), .A2(execstage_BusA[6]), .B1(n16356), .B2(n2814), 
        .ZN(n2786) );
  XOR2_X2 U8096 ( .A(n13116), .B(n6028), .Z(n2814) );
  AOI22_X2 U8098 ( .A1(n6030), .A2(execstage_BusA[5]), .B1(n2836), .B2(n2837), 
        .ZN(n2813) );
  XOR2_X2 U8099 ( .A(n13119), .B(n6030), .Z(n2837) );
  OAI22_X2 U8100 ( .A1(n16450), .A2(n8738), .B1(n2859), .B2(n2858), .ZN(n2836)
         );
  XOR2_X2 U8101 ( .A(n8738), .B(n6032), .Z(n2858) );
  AOI22_X2 U8102 ( .A1(n6033), .A2(n8651), .B1(n16479), .B2(n2890), .ZN(n2859)
         );
  XOR2_X2 U8103 ( .A(n8651), .B(n6033), .Z(n2890) );
  AOI22_X2 U8105 ( .A1(n6035), .A2(execstage_BusA[2]), .B1(n3417), .B2(n3416), 
        .ZN(n6034) );
  XOR2_X2 U8106 ( .A(execstage_BusA[2]), .B(n6035), .Z(n3416) );
  OAI22_X2 U8107 ( .A1(n6036), .A2(n13151), .B1(n4940), .B2(n4939), .ZN(n3417)
         );
  XOR2_X2 U8108 ( .A(n6036), .B(execstage_BusA[1]), .Z(n4939) );
  AOI22_X2 U8109 ( .A1(n6037), .A2(n13795), .B1(n6038), .B2(execstage_ALU_sel), 
        .ZN(n4940) );
  XOR2_X2 U8110 ( .A(n13132), .B(n13197), .Z(n6036) );
  XOR2_X2 U8111 ( .A(n13132), .B(n13174), .Z(n6035) );
  XNOR2_X2 U8112 ( .A(n13134), .B(n13203), .ZN(n6033) );
  XNOR2_X2 U8114 ( .A(n13134), .B(n13192), .ZN(n6032) );
  XOR2_X2 U8115 ( .A(n13132), .B(n13205), .Z(n6030) );
  XNOR2_X2 U8116 ( .A(n13134), .B(n13211), .ZN(n6028) );
  XOR2_X2 U8117 ( .A(n13132), .B(n13214), .Z(n6027) );
  XOR2_X2 U8118 ( .A(n13132), .B(n13215), .Z(n6026) );
  XNOR2_X2 U8119 ( .A(n13134), .B(n13158), .ZN(n6024) );
  XOR2_X2 U8120 ( .A(n13135), .B(n5800), .Z(n5799) );
  XNOR2_X2 U8121 ( .A(n13134), .B(n13161), .ZN(n5800) );
  AOI221_X2 U8124 ( .B1(n6042), .B2(n13783), .C1(n8807), .C2(n13129), .A(n6043), .ZN(n6041) );
  OAI22_X2 U8125 ( .A1(n2896), .A2(n5619), .B1(n2721), .B2(n6044), .ZN(n6043)
         );
  NAND2_X2 U8126 ( .A1(n6045), .A2(execstage_AluCtrl[1]), .ZN(n2721) );
  NAND2_X2 U8133 ( .A1(n21), .A2(n6049), .ZN(execstage_ALU_N160) );
  NAND4_X2 U8134 ( .A1(execstage_AluCtrl[0]), .A2(execstage_AluCtrl[1]), .A3(
        n8697), .A4(n8660), .ZN(n6049) );
  NAND2_X2 U8135 ( .A1(n6051), .A2(n8660), .ZN(n21) );
  XOR2_X2 U8136 ( .A(execstage_ALU_sel), .B(n6038), .Z(n6042) );
  XOR2_X2 U8137 ( .A(n13795), .B(n6037), .Z(n6038) );
  XNOR2_X2 U8138 ( .A(n13132), .B(n13129), .ZN(n6037) );
  AOI221_X2 U8140 ( .B1(n13105), .B2(n4388), .C1(n6052), .C2(n6053), .A(n6054), 
        .ZN(n6040) );
  NOR4_X2 U8141 ( .A1(execstage_AluCtrl[3]), .A2(n6055), .A3(n8697), .A4(n8720), .ZN(n6054) );
  NOR4_X2 U8150 ( .A1(n6066), .A2(n2902), .A3(n5796), .A4(n16533), .ZN(n6065)
         );
  NAND2_X2 U8152 ( .A1(n6068), .A2(n5619), .ZN(n6044) );
  NAND2_X2 U8153 ( .A1(n13795), .A2(n13129), .ZN(n5619) );
  NAND4_X2 U8154 ( .A1(n6069), .A2(n5535), .A3(n6070), .A4(n5717), .ZN(n6066)
         );
  XNOR2_X2 U8158 ( .A(n6077), .B(n2902), .ZN(n6062) );
  OAI22_X2 U8159 ( .A1(execstage_ALU_ra_row2_31_), .A2(n6078), .B1(n6079), 
        .B2(n2902), .ZN(n6077) );
  AOI22_X2 U8160 ( .A1(n16436), .A2(n6081), .B1(n16437), .B2(n8658), .ZN(n6079) );
  OAI221_X2 U8161 ( .B1(n6082), .B2(n16421), .C1(execstage_BusA[29]), .C2(
        n2970), .A(n6084), .ZN(n6081) );
  OR3_X2 U8165 ( .A1(n2946), .A2(execstage_BusA[26]), .A3(n3953), .ZN(n6088)
         );
  AOI22_X2 U8166 ( .A1(n16434), .A2(n6090), .B1(n16435), .B2(n8732), .ZN(n6082) );
  OAI22_X2 U8167 ( .A1(execstage_BusA[24]), .A2(n3480), .B1(n6091), .B2(n4394), 
        .ZN(n6090) );
  AOI22_X2 U8168 ( .A1(n16430), .A2(n6093), .B1(n16431), .B2(n8656), .ZN(n6091) );
  OAI211_X2 U8169 ( .C1(n6094), .C2(n6074), .A(n6095), .B(n6096), .ZN(n6093)
         );
  AOI22_X2 U8170 ( .A1(n16411), .A2(n6098), .B1(n13111), .B2(n8653), .ZN(n6096) );
  OAI22_X2 U8171 ( .A1(execstage_BusA[21]), .A2(n3500), .B1(n6099), .B2(n4799), 
        .ZN(n6098) );
  AOI22_X2 U8172 ( .A1(n16408), .A2(n6101), .B1(n16409), .B2(n13117), .ZN(
        n6099) );
  OR3_X2 U8174 ( .A1(n13110), .A2(execstage_BusA[18]), .A3(n5058), .ZN(n6102)
         );
  AOI22_X2 U8176 ( .A1(n16419), .A2(n6105), .B1(n13107), .B2(n8734), .ZN(n6094) );
  OAI22_X2 U8177 ( .A1(execstage_BusA[15]), .A2(n13167), .B1(n16359), .B2(
        n6106), .ZN(n6105) );
  AOI22_X2 U8178 ( .A1(n6107), .A2(n5535), .B1(n13179), .B2(n8657), .ZN(n6106)
         );
  OAI22_X2 U8179 ( .A1(n8655), .A2(n13165), .B1(n16364), .B2(n6108), .ZN(n6107) );
  AOI22_X2 U8180 ( .A1(n6109), .A2(n5717), .B1(n13164), .B2(n8695), .ZN(n6108)
         );
  OAI22_X2 U8181 ( .A1(n13121), .A2(n13180), .B1(n5796), .B2(n6110), .ZN(n6109) );
  AOI221_X2 U8182 ( .B1(n13161), .B2(n13136), .C1(n6076), .C2(n6111), .A(n6112), .ZN(n6110) );
  OAI221_X2 U8184 ( .B1(n6113), .B2(n6072), .C1(execstage_BusA[8]), .C2(n13215), .A(n6114), .ZN(n6111) );
  AOI22_X2 U8185 ( .A1(n6115), .A2(n6116), .B1(n6117), .B2(n16329), .ZN(n6114)
         );
  OAI22_X2 U8186 ( .A1(execstage_BusA[7]), .A2(n13212), .B1(n2791), .B2(n6119), 
        .ZN(n6117) );
  AOI22_X2 U8187 ( .A1(n6120), .A2(n16413), .B1(n13211), .B2(n13154), .ZN(
        n6119) );
  AOI221_X2 U8192 ( .B1(n13177), .B2(n13793), .C1(n6124), .C2(n13129), .A(
        n6125), .ZN(n6113) );
  XNOR2_X2 U8194 ( .A(n6126), .B(n2902), .ZN(n6059) );
  OAI22_X2 U8195 ( .A1(n16438), .A2(n8744), .B1(n6127), .B2(n2902), .ZN(n6126)
         );
  XOR2_X2 U8196 ( .A(n8744), .B(n6078), .Z(n2902) );
  OAI221_X2 U8198 ( .B1(n6132), .B2(n6074), .C1(n13111), .C2(n8653), .A(n6133), 
        .ZN(n6131) );
  OAI22_X2 U8202 ( .A1(n16406), .A2(n8646), .B1(n6137), .B2(n4799), .ZN(n6134)
         );
  AOI22_X2 U8203 ( .A1(n16408), .A2(n6138), .B1(execstage_BusA[20]), .B2(n3178), .ZN(n6137) );
  OAI22_X2 U8204 ( .A1(n13112), .A2(n8654), .B1(n5058), .B2(n6139), .ZN(n6138)
         );
  NAND2_X2 U8205 ( .A1(execstage_BusA[18]), .A2(n13110), .ZN(n6139) );
  OR2_X2 U8210 ( .A1(n16388), .A2(n5268), .ZN(n6074) );
  XOR2_X2 U8211 ( .A(n8647), .B(n3529), .Z(n5268) );
  NOR4_X2 U8215 ( .A1(n5163), .A2(n4673), .A3(n6141), .A4(n4799), .ZN(n6103)
         );
  XOR2_X2 U8216 ( .A(n8646), .B(n3500), .Z(n4799) );
  OR2_X2 U8219 ( .A1(n5058), .A2(n4917), .ZN(n6141) );
  XNOR2_X2 U8220 ( .A(n13117), .B(n16409), .ZN(n4917) );
  XOR2_X2 U8223 ( .A(n8654), .B(n3515), .Z(n5058) );
  XNOR2_X2 U8226 ( .A(n8653), .B(n13111), .ZN(n4673) );
  XOR2_X2 U8229 ( .A(n8650), .B(n3201), .Z(n5163) );
  AOI22_X2 U8231 ( .A1(n16419), .A2(n6142), .B1(execstage_BusA[16]), .B2(
        n13108), .ZN(n6132) );
  OAI22_X2 U8232 ( .A1(n13168), .A2(n8645), .B1(n16359), .B2(n6143), .ZN(n6142) );
  AOI22_X2 U8233 ( .A1(n6144), .A2(n5535), .B1(execstage_BusA[14]), .B2(n13178), .ZN(n6143) );
  NAND2_X2 U8234 ( .A1(n5526), .A2(n3625), .ZN(n5535) );
  NAND2_X2 U8235 ( .A1(n13179), .A2(execstage_BusA[14]), .ZN(n3625) );
  NAND2_X2 U8237 ( .A1(n8657), .A2(n13178), .ZN(n5526) );
  OAI22_X2 U8238 ( .A1(execstage_Imm32[14]), .A2(n13785), .B1(n13788), .B2(
        busB_1[14]), .ZN(n3293) );
  OAI22_X2 U8239 ( .A1(n13166), .A2(n8710), .B1(n16364), .B2(n6145), .ZN(n6144) );
  AOI22_X2 U8240 ( .A1(n6146), .A2(n5717), .B1(execstage_BusA[12]), .B2(n13162), .ZN(n6145) );
  NAND2_X2 U8241 ( .A1(n5648), .A2(n4237), .ZN(n5717) );
  NAND2_X2 U8242 ( .A1(n13164), .A2(execstage_BusA[12]), .ZN(n4237) );
  NAND2_X2 U8244 ( .A1(n8695), .A2(n13162), .ZN(n5648) );
  OAI22_X2 U8245 ( .A1(execstage_Imm32[12]), .A2(n13785), .B1(execstage_ALUSrc), .B2(busB_1[12]), .ZN(n3555) );
  OAI22_X2 U8246 ( .A1(n13182), .A2(n8736), .B1(n5796), .B2(n6147), .ZN(n6146)
         );
  AOI221_X2 U8247 ( .B1(n13122), .B2(n13159), .C1(n6076), .C2(n6148), .A(n6149), .ZN(n6147) );
  OAI221_X2 U8249 ( .B1(n6150), .B2(n6072), .C1(n13217), .C2(n13148), .A(n6151), .ZN(n6148) );
  AND3_X2 U8251 ( .A1(n6116), .A2(n13201), .A3(n13791), .ZN(n6153) );
  OAI22_X2 U8253 ( .A1(n13214), .A2(n13155), .B1(n2791), .B2(n6154), .ZN(n6152) );
  AOI22_X2 U8254 ( .A1(n6155), .A2(n16413), .B1(execstage_BusA[6]), .B2(n13209), .ZN(n6154) );
  NAND2_X2 U8261 ( .A1(n6116), .A2(n2895), .ZN(n6072) );
  NAND2_X2 U8262 ( .A1(n2887), .A2(n2897), .ZN(n2895) );
  NAND2_X2 U8263 ( .A1(n13204), .A2(n13791), .ZN(n2897) );
  NAND2_X2 U8264 ( .A1(n13790), .A2(n13201), .ZN(n2887) );
  OR3_X2 U8267 ( .A1(n2791), .A2(n2840), .A3(n2817), .ZN(n6157) );
  NAND2_X2 U8270 ( .A1(n13211), .A2(n13116), .ZN(n5606) );
  OAI22_X2 U8273 ( .A1(execstage_Imm32[6]), .A2(n13785), .B1(execstage_ALUSrc), 
        .B2(busB_1[6]), .ZN(n2804) );
  NAND2_X2 U8276 ( .A1(n13207), .A2(n13119), .ZN(n5778) );
  OAI22_X2 U8279 ( .A1(execstage_Imm32[5]), .A2(n13785), .B1(execstage_ALUSrc), 
        .B2(busB_1[5]), .ZN(n2830) );
  NAND2_X2 U8282 ( .A1(n13214), .A2(execstage_BusA[7]), .ZN(n5440) );
  OAI22_X2 U8285 ( .A1(execstage_Imm32[7]), .A2(n13785), .B1(execstage_ALUSrc), 
        .B2(busB_1[7]), .ZN(n2775) );
  NAND2_X2 U8288 ( .A1(n13217), .A2(execstage_BusA[8]), .ZN(n5259) );
  OAI22_X2 U8291 ( .A1(execstage_Imm32[8]), .A2(n13786), .B1(execstage_ALUSrc), 
        .B2(busB_1[8]), .ZN(n2748) );
  NAND2_X2 U8292 ( .A1(n8738), .A2(n13190), .ZN(n2849) );
  NAND2_X2 U8294 ( .A1(execstage_BusA[4]), .A2(n13192), .ZN(n2861) );
  AND2_X2 U8299 ( .A1(n4925), .A2(n6010), .ZN(n4947) );
  NAND2_X2 U8300 ( .A1(n13198), .A2(execstage_BusA[1]), .ZN(n6010) );
  NAND2_X2 U8301 ( .A1(n13151), .A2(n13196), .ZN(n4925) );
  NAND2_X2 U8308 ( .A1(n13161), .A2(n13122), .ZN(n4790) );
  NAND2_X2 U8313 ( .A1(n13158), .A2(n8648), .ZN(n5048) );
  OAI22_X2 U8315 ( .A1(execstage_Imm32[9]), .A2(n13786), .B1(execstage_ALUSrc), 
        .B2(busB_1[9]), .ZN(n3569) );
  OAI22_X2 U8317 ( .A1(execstage_Imm32[10]), .A2(n13786), .B1(execstage_ALUSrc), .B2(busB_1[10]), .ZN(n3565) );
  NAND2_X2 U8320 ( .A1(n13182), .A2(n13121), .ZN(n4522) );
  OAI22_X2 U8324 ( .A1(execstage_Imm32[11]), .A2(n13786), .B1(execstage_ALUSrc), .B2(busB_1[11]), .ZN(n3130) );
  NAND2_X2 U8326 ( .A1(n5609), .A2(n3939), .ZN(n6070) );
  NAND2_X2 U8327 ( .A1(n13166), .A2(n8655), .ZN(n3939) );
  NAND2_X2 U8328 ( .A1(n8710), .A2(n13165), .ZN(n5609) );
  OAI22_X2 U8331 ( .A1(execstage_Imm32[13]), .A2(n13786), .B1(execstage_ALUSrc), .B2(busB_1[13]), .ZN(n3548) );
  NAND2_X2 U8333 ( .A1(n5442), .A2(n3196), .ZN(n6069) );
  NAND2_X2 U8334 ( .A1(n13168), .A2(execstage_BusA[15]), .ZN(n3196) );
  NAND2_X2 U8335 ( .A1(n8645), .A2(n13167), .ZN(n5442) );
  OAI22_X2 U8338 ( .A1(execstage_Imm32[15]), .A2(n13786), .B1(execstage_ALUSrc), .B2(busB_1[15]), .ZN(n3543) );
  XNOR2_X2 U8340 ( .A(n13139), .B(n13107), .ZN(n5360) );
  NAND4_X2 U8344 ( .A1(n16436), .A2(n6160), .A3(n6161), .A4(n16430), .ZN(n6073) );
  XNOR2_X2 U8346 ( .A(n8656), .B(n16431), .ZN(n4533) );
  OAI221_X2 U8350 ( .B1(n6162), .B2(n16421), .C1(n16424), .C2(n8737), .A(n6163), .ZN(n6129) );
  OAI22_X2 U8354 ( .A1(n16427), .A2(n8713), .B1(n3953), .B2(n6166), .ZN(n6164)
         );
  NAND2_X2 U8355 ( .A1(execstage_BusA[26]), .A2(n2946), .ZN(n6166) );
  XNOR2_X2 U8361 ( .A(n8737), .B(n16424), .ZN(n3442) );
  OAI22_X2 U8363 ( .A1(execstage_Imm32[29]), .A2(n13786), .B1(n13788), .B2(
        busB_1[29]), .ZN(n2970) );
  XOR2_X2 U8364 ( .A(n8735), .B(n3455), .Z(n3632) );
  OAI22_X2 U8365 ( .A1(execstage_Imm32[28]), .A2(n13786), .B1(execstage_ALUSrc), .B2(busB_1[28]), .ZN(n3455) );
  XOR2_X2 U8367 ( .A(n8713), .B(n3209), .Z(n3953) );
  OAI22_X2 U8368 ( .A1(execstage_Imm32[27]), .A2(n13786), .B1(n13788), .B2(
        busB_1[27]), .ZN(n3209) );
  XOR2_X2 U8370 ( .A(n8733), .B(n2946), .Z(n4105) );
  AOI22_X2 U8373 ( .A1(n16434), .A2(n6168), .B1(execstage_BusA[25]), .B2(n3474), .ZN(n6162) );
  OAI22_X2 U8374 ( .A1(n16433), .A2(n8731), .B1(n4394), .B2(n6169), .ZN(n6168)
         );
  NAND2_X2 U8375 ( .A1(execstage_BusA[23]), .A2(n3004), .ZN(n6169) );
  XOR2_X2 U8377 ( .A(execstage_BusA[24]), .B(n16433), .Z(n4394) );
  XNOR2_X2 U8382 ( .A(n8732), .B(n16435), .ZN(n4248) );
  OAI22_X2 U8384 ( .A1(execstage_Imm32[25]), .A2(n13787), .B1(n13788), .B2(
        busB_1[25]), .ZN(n3474) );
  XNOR2_X2 U8387 ( .A(n8658), .B(n16437), .ZN(n3227) );
  OAI22_X2 U8389 ( .A1(execstage_Imm32[30]), .A2(n13787), .B1(n13788), .B2(
        busB_1[30]), .ZN(n6128) );
  OAI22_X2 U8392 ( .A1(execstage_Imm32[31]), .A2(n13787), .B1(n13788), .B2(
        busB_1[31]), .ZN(n6078) );
  NAND2_X2 U8394 ( .A1(n16549), .A2(n13190), .ZN(n5642) );
  NAND2_X2 U8396 ( .A1(execstage_AluCtrl[3]), .A2(n6051), .ZN(n3429) );
  AOI22_X2 U8398 ( .A1(n13218), .A2(n6068), .B1(n6170), .B2(n3403), .ZN(n6039)
         );
  NAND2_X2 U8399 ( .A1(n3653), .A2(n3222), .ZN(n3403) );
  OR4_X2 U8400 ( .A1(n8660), .A2(n8720), .A3(n8697), .A4(execstage_AluCtrl[0]), 
        .ZN(n3222) );
  NAND2_X2 U8401 ( .A1(n6047), .A2(execstage_AluCtrl[3]), .ZN(n3653) );
  AND3_X2 U8402 ( .A1(execstage_AluCtrl[2]), .A2(n8720), .A3(
        execstage_AluCtrl[0]), .ZN(n6047) );
  OAI222_X2 U8403 ( .A1(n6171), .A2(n3231), .B1(n13192), .B2(n6172), .C1(
        n16401), .C2(n2909), .ZN(n6170) );
  OAI221_X2 U8405 ( .B1(n16507), .B2(n13104), .C1(n16506), .C2(n5160), .A(
        n6175), .ZN(n5359) );
  AOI22_X2 U8406 ( .A1(n8659), .A2(n2749), .B1(n16471), .B2(n2753), .ZN(n6175)
         );
  OAI221_X2 U8407 ( .B1(n13186), .B2(n8653), .C1(n13169), .C2(n8730), .A(n6176), .ZN(n2753) );
  NAND2_X2 U8410 ( .A1(n16534), .A2(n13199), .ZN(n4101) );
  NAND2_X2 U8412 ( .A1(execstage_BusA[23]), .A2(n13129), .ZN(n4490) );
  NAND2_X2 U8414 ( .A1(execstage_BusA[21]), .A2(n13129), .ZN(n4764) );
  OAI221_X2 U8417 ( .B1(n13186), .B2(n8650), .C1(n8734), .C2(n3434), .A(n6177), 
        .ZN(n2749) );
  AOI22_X2 U8418 ( .A1(n16404), .A2(n13198), .B1(n16536), .B2(n13195), .ZN(
        n6177) );
  NAND2_X2 U8420 ( .A1(execstage_BusA[17]), .A2(n13129), .ZN(n5131) );
  NAND2_X2 U8422 ( .A1(execstage_BusA[19]), .A2(n13102), .ZN(n4884) );
  OAI211_X2 U8426 ( .C1(n13185), .C2(n8658), .A(n6178), .B(n6179), .ZN(n3652)
         );
  AOI22_X2 U8427 ( .A1(n3238), .A2(n13195), .B1(execstage_BusA[28]), .B2(
        n13171), .ZN(n6179) );
  NAND2_X2 U8436 ( .A1(n16537), .A2(n13199), .ZN(n3242) );
  NAND2_X2 U8438 ( .A1(execstage_BusA[27]), .A2(n13102), .ZN(n3641) );
  NAND2_X2 U8440 ( .A1(execstage_BusA[25]), .A2(n13129), .ZN(n4205) );
  NAND2_X2 U8441 ( .A1(execstage_BusA[26]), .A2(n13183), .ZN(n3640) );
  NAND2_X2 U8442 ( .A1(execstage_BusA[24]), .A2(n13171), .ZN(n4389) );
  OAI211_X2 U8444 ( .C1(n13194), .C2(n3412), .A(n5644), .B(n6181), .ZN(n2854)
         );
  AOI22_X2 U8445 ( .A1(n16539), .A2(n13195), .B1(n13187), .B2(
        execstage_BusA[6]), .ZN(n6181) );
  NAND2_X2 U8447 ( .A1(execstage_BusA[5]), .A2(n13102), .ZN(n3408) );
  NAND2_X2 U8448 ( .A1(n13171), .A2(execstage_BusA[4]), .ZN(n5644) );
  NAND2_X2 U8450 ( .A1(n13115), .A2(n13102), .ZN(n3412) );
  OAI221_X2 U8453 ( .B1(n13136), .B2(n13184), .C1(n13148), .C2(n13170), .A(
        n6182), .ZN(n2750) );
  AOI22_X2 U8454 ( .A1(n16542), .A2(n13198), .B1(n16541), .B2(n13195), .ZN(
        n6182) );
  NAND2_X2 U8456 ( .A1(n13118), .A2(n13102), .ZN(n3411) );
  NAND2_X2 U8458 ( .A1(n13121), .A2(n13102), .ZN(n5692) );
  OAI221_X2 U8463 ( .B1(n13138), .B2(n13184), .C1(n8695), .C2(n3434), .A(n6183), .ZN(n2751) );
  AOI22_X2 U8464 ( .A1(n16544), .A2(n13198), .B1(n16543), .B2(n13195), .ZN(
        n6183) );
  NAND2_X2 U8466 ( .A1(n13120), .A2(n13102), .ZN(n5505) );
  NAND2_X2 U8468 ( .A1(execstage_BusA[15]), .A2(n13102), .ZN(n5326) );
  NAND2_X2 U8472 ( .A1(n13204), .A2(n13177), .ZN(n5160) );
  NAND2_X2 U8476 ( .A1(n8659), .A2(n2909), .ZN(n3231) );
  OAI22_X2 U8477 ( .A1(execstage_Imm32[4]), .A2(n13787), .B1(n13788), .B2(
        busB_1[4]), .ZN(n2909) );
  OAI22_X2 U8480 ( .A1(execstage_Imm32[3]), .A2(n13787), .B1(n13788), .B2(
        busB_1[3]), .ZN(n2869) );
  OAI22_X2 U8481 ( .A1(execstage_Imm32[2]), .A2(n13787), .B1(n13788), .B2(
        busB_1[2]), .ZN(n3338) );
  NOR4_X2 U8482 ( .A1(n16516), .A2(n4388), .A3(n6009), .A4(n16512), .ZN(n6171)
         );
  NAND2_X2 U8484 ( .A1(n13187), .A2(n13792), .ZN(n5643) );
  NAND2_X2 U8486 ( .A1(n13198), .A2(n5264), .ZN(n2919) );
  NAND2_X2 U8489 ( .A1(n13791), .A2(n13102), .ZN(n5646) );
  NAND2_X2 U8492 ( .A1(n13196), .A2(n5264), .ZN(n3434) );
  NAND2_X2 U8494 ( .A1(n4928), .A2(n13196), .ZN(n6020) );
  OAI22_X2 U8495 ( .A1(execstage_Imm32[1]), .A2(n13787), .B1(n13788), .B2(
        busB_1[1]), .ZN(n2881) );
  NAND2_X2 U8498 ( .A1(n8712), .A2(n5264), .ZN(n6068) );
  NAND2_X2 U8509 ( .A1(N43), .A2(N27), .ZN(N47) );
  AND3_X2 U8510 ( .A1(N34), .A2(n6186), .A3(regwrite_2), .ZN(N44) );
  NAND2_X2 U8511 ( .A1(N38), .A2(n16215), .ZN(N43) );
  NAND2_X2 U8513 ( .A1(regwrite_1), .A2(N32), .ZN(n6186) );
  AND3_X2 U8514 ( .A1(regwrite_2), .A2(n6187), .A3(N19), .ZN(N28) );
  NAND2_X2 U8515 ( .A1(N23), .A2(n16216), .ZN(N27) );
  NAND2_X2 U8517 ( .A1(N17), .A2(regwrite_1), .ZN(n6187) );
  OAI22_X2 U8518 ( .A1(n13809), .A2(n6188), .B1(N15), .B2(n16371), .ZN(N14) );
  INV_X4 U8520 ( .A(N15), .ZN(n6188) );
  NAND4_X2 U8523 ( .A1(instruction_2[29]), .A2(instruction_2[28]), .A3(n6191), 
        .A4(instruction_2[27]), .ZN(n6190) );
  AND2_X4 U8529 ( .A1(n6047), .A2(n8660), .ZN(n8649) );
  AND2_X4 U8530 ( .A1(n13174), .A2(n13201), .ZN(n8659) );
  AND2_X4 U8531 ( .A1(n664), .A2(n495), .ZN(n8661) );
  AND2_X4 U8532 ( .A1(n836), .A2(n495), .ZN(n8662) );
  AND2_X4 U8533 ( .A1(n836), .A2(n564), .ZN(n8663) );
  AND2_X4 U8534 ( .A1(n836), .A2(n529), .ZN(n8664) );
  AND2_X4 U8535 ( .A1(n664), .A2(n564), .ZN(n8665) );
  AND2_X4 U8536 ( .A1(n664), .A2(n529), .ZN(n8666) );
  AND2_X4 U8537 ( .A1(n530), .A2(n495), .ZN(n8667) );
  AND2_X4 U8538 ( .A1(n1571), .A2(n733), .ZN(n8668) );
  AND2_X4 U8539 ( .A1(n1571), .A2(n699), .ZN(n8669) );
  AND2_X4 U8540 ( .A1(n2407), .A2(n733), .ZN(n8670) );
  AND2_X4 U8541 ( .A1(n2407), .A2(n699), .ZN(n8671) );
  AND2_X4 U8542 ( .A1(n2273), .A2(n733), .ZN(n8672) );
  AND2_X4 U8543 ( .A1(n2273), .A2(n699), .ZN(n8673) );
  AND2_X4 U8544 ( .A1(n2106), .A2(n733), .ZN(n8674) );
  AND2_X4 U8545 ( .A1(n2106), .A2(n699), .ZN(n8675) );
  AND2_X4 U8546 ( .A1(n1973), .A2(n733), .ZN(n8676) );
  AND2_X4 U8547 ( .A1(n1973), .A2(n699), .ZN(n8677) );
  AND2_X4 U8548 ( .A1(n1772), .A2(n733), .ZN(n8678) );
  AND2_X4 U8549 ( .A1(n1806), .A2(n733), .ZN(n8679) );
  AND2_X4 U8550 ( .A1(n1806), .A2(n699), .ZN(n8680) );
  AND2_X4 U8551 ( .A1(n1772), .A2(n699), .ZN(n8681) );
  AND2_X4 U8552 ( .A1(n1638), .A2(n733), .ZN(n8682) );
  AND2_X4 U8553 ( .A1(n1638), .A2(n699), .ZN(n8683) );
  AND2_X4 U8554 ( .A1(n1169), .A2(n733), .ZN(n8684) );
  AND2_X4 U8555 ( .A1(n1169), .A2(n699), .ZN(n8685) );
  AND2_X4 U8556 ( .A1(n1003), .A2(n733), .ZN(n8686) );
  AND2_X4 U8557 ( .A1(n1003), .A2(n699), .ZN(n8687) );
  AND2_X4 U8558 ( .A1(n870), .A2(n733), .ZN(n8688) );
  AND2_X4 U8559 ( .A1(n870), .A2(n699), .ZN(n8689) );
  AND2_X4 U8560 ( .A1(n698), .A2(n733), .ZN(n8690) );
  AND2_X4 U8561 ( .A1(n698), .A2(n699), .ZN(n8691) );
  AND2_X4 U8562 ( .A1(n13204), .A2(n13174), .ZN(n8696) );
  AND2_X4 U8563 ( .A1(n836), .A2(n460), .ZN(n8698) );
  AND2_X4 U8564 ( .A1(n664), .A2(n460), .ZN(n8699) );
  AND2_X4 U8565 ( .A1(n530), .A2(n460), .ZN(n8700) );
  AND2_X4 U8566 ( .A1(n564), .A2(n461), .ZN(n8701) );
  AND2_X4 U8567 ( .A1(n529), .A2(n461), .ZN(n8702) );
  AND2_X4 U8568 ( .A1(n564), .A2(n530), .ZN(n8703) );
  AND2_X4 U8569 ( .A1(n529), .A2(n530), .ZN(n8704) );
  AND2_X4 U8570 ( .A1(n495), .A2(n461), .ZN(n8705) );
  AND2_X4 U8571 ( .A1(n460), .A2(n461), .ZN(n8706) );
  OR2_X4 U8572 ( .A1(n3653), .A2(n2909), .ZN(n8722) );
  INV_X4 U8573 ( .A(n10943), .ZN(n10947) );
  INV_X4 U8574 ( .A(n10943), .ZN(n10950) );
  INV_X4 U8575 ( .A(n10943), .ZN(n10944) );
  INV_X4 U8576 ( .A(n10943), .ZN(n10951) );
  INV_X4 U8577 ( .A(n10943), .ZN(n10945) );
  INV_X4 U8578 ( .A(n10943), .ZN(n10948) );
  INV_X4 U8579 ( .A(n10943), .ZN(n10949) );
  INV_X4 U8580 ( .A(n10943), .ZN(n10946) );
  OAI21_X2 U8581 ( .B1(n4603), .B2(n4604), .A(n4524), .ZN(n4602) );
  INV_X4 U8582 ( .A(n13095), .ZN(n13086) );
  INV_X4 U8583 ( .A(n13095), .ZN(n13091) );
  INV_X4 U8584 ( .A(n13095), .ZN(n13085) );
  INV_X4 U8585 ( .A(n13095), .ZN(n13090) );
  INV_X4 U8586 ( .A(n13095), .ZN(n13084) );
  INV_X4 U8587 ( .A(n13095), .ZN(n13089) );
  INV_X4 U8588 ( .A(n13095), .ZN(n13088) );
  INV_X4 U8589 ( .A(n13095), .ZN(n13087) );
  INV_X4 U8590 ( .A(n2785), .ZN(n16455) );
  INV_X4 U8591 ( .A(n4929), .ZN(n16449) );
  INV_X4 U8592 ( .A(n2772), .ZN(n16448) );
  INV_X4 U8593 ( .A(decode_rs2_3_), .ZN(n10943) );
  INV_X4 U8594 ( .A(n10955), .ZN(n10957) );
  INV_X4 U8595 ( .A(n10955), .ZN(n10960) );
  INV_X4 U8596 ( .A(n10955), .ZN(n10958) );
  INV_X4 U8597 ( .A(n10955), .ZN(n10959) );
  INV_X4 U8598 ( .A(n10955), .ZN(n10956) );
  INV_X4 U8599 ( .A(n10943), .ZN(n10953) );
  INV_X4 U8600 ( .A(n10943), .ZN(n10954) );
  INV_X4 U8601 ( .A(n10943), .ZN(n10952) );
  AOI21_X2 U8602 ( .B1(n5837), .B2(n5838), .A(n5841), .ZN(n5751) );
  AOI21_X2 U8603 ( .B1(n4965), .B2(n4966), .A(n4967), .ZN(n4826) );
  AOI21_X2 U8604 ( .B1(n4693), .B2(n4694), .A(n4695), .ZN(n4562) );
  OAI21_X2 U8605 ( .B1(n13189), .B2(n13154), .A(n5890), .ZN(n5889) );
  OAI21_X2 U8606 ( .B1(n13189), .B2(n13135), .A(n5498), .ZN(n5497) );
  OAI21_X2 U8607 ( .B1(n5734), .B2(n5735), .A(n5706), .ZN(n5733) );
  OAI21_X2 U8608 ( .B1(n5375), .B2(n5376), .A(n5351), .ZN(n5374) );
  OAI21_X2 U8609 ( .B1(n5935), .B2(n5936), .A(n5937), .ZN(n5934) );
  OAI21_X2 U8610 ( .B1(n5886), .B2(n5885), .A(n5938), .ZN(n5884) );
  OAI21_X2 U8611 ( .B1(n16315), .B2(n5396), .A(n5397), .ZN(n5304) );
  OAI21_X2 U8612 ( .B1(n5294), .B2(n5295), .A(n5296), .ZN(n5200) );
  OAI21_X2 U8613 ( .B1(n3878), .B2(n3879), .A(n3880), .ZN(n3729) );
  OAI21_X2 U8614 ( .B1(n16268), .B2(n4167), .A(n4168), .ZN(n4018) );
  OAI21_X2 U8615 ( .B1(n16267), .B2(n4162), .A(n4163), .ZN(n4013) );
  OAI21_X2 U8616 ( .B1(n3865), .B2(n3866), .A(n3867), .ZN(n3714) );
  OAI21_X2 U8617 ( .B1(n5390), .B2(n5391), .A(n5392), .ZN(n5299) );
  OAI21_X2 U8618 ( .B1(n16271), .B2(n4034), .A(n4035), .ZN(n3883) );
  OAI21_X2 U8619 ( .B1(n5289), .B2(n5290), .A(n5291), .ZN(n5195) );
  OAI21_X2 U8620 ( .B1(n5424), .B2(n5425), .A(n5426), .ZN(n5329) );
  OAI21_X2 U8621 ( .B1(n5771), .B2(n5772), .A(n5773), .ZN(n5695) );
  OAI21_X2 U8622 ( .B1(n5774), .B2(n5775), .A(n5776), .ZN(n5698) );
  OAI21_X2 U8623 ( .B1(n5599), .B2(n5600), .A(n5601), .ZN(n5514) );
  OAI21_X2 U8624 ( .B1(n5427), .B2(n5428), .A(n5429), .ZN(n5332) );
  OAI21_X2 U8625 ( .B1(n5602), .B2(n5603), .A(n5604), .ZN(n5517) );
  OAI21_X2 U8626 ( .B1(n5430), .B2(n5431), .A(n5432), .ZN(n5335) );
  OAI21_X2 U8627 ( .B1(n5246), .B2(n5247), .A(n5248), .ZN(n5140) );
  OAI21_X2 U8628 ( .B1(n5249), .B2(n5250), .A(n5251), .ZN(n5143) );
  OAI21_X2 U8629 ( .B1(n5033), .B2(n5034), .A(n5035), .ZN(n4893) );
  OAI21_X2 U8630 ( .B1(n5252), .B2(n5253), .A(n5254), .ZN(n5146) );
  OAI21_X2 U8631 ( .B1(n16338), .B2(n5256), .A(n5257), .ZN(n5149) );
  OAI21_X2 U8632 ( .B1(n5039), .B2(n5040), .A(n5041), .ZN(n4899) );
  OAI21_X2 U8633 ( .B1(n5042), .B2(n5043), .A(n5044), .ZN(n4902) );
  OAI21_X2 U8634 ( .B1(n4778), .B2(n4779), .A(n4780), .ZN(n4646) );
  OAI21_X2 U8635 ( .B1(n5045), .B2(n5046), .A(n5047), .ZN(n4905) );
  OAI21_X2 U8636 ( .B1(n4784), .B2(n4785), .A(n4786), .ZN(n4652) );
  OAI21_X2 U8637 ( .B1(n4787), .B2(n4788), .A(n4789), .ZN(n4655) );
  OAI21_X2 U8638 ( .B1(n4513), .B2(n4514), .A(n4515), .ZN(n4374) );
  OAI21_X2 U8639 ( .B1(n4519), .B2(n4520), .A(n4521), .ZN(n4380) );
  OAI21_X2 U8640 ( .B1(n16475), .B2(n5594), .A(n5595), .ZN(n5508) );
  OAI21_X2 U8641 ( .B1(n5436), .B2(n5437), .A(n5438), .ZN(n5341) );
  OAI21_X2 U8642 ( .B1(n4231), .B2(n4232), .A(n4233), .ZN(n4089) );
  OAI21_X2 U8643 ( .B1(n3253), .B2(n3254), .A(n2949), .ZN(n2963) );
  OAI21_X2 U8644 ( .B1(n5887), .B2(n5888), .A(n5926), .ZN(n5875) );
  OAI21_X2 U8645 ( .B1(n16344), .B2(n5846), .A(n5866), .ZN(n5864) );
  OAI21_X2 U8646 ( .B1(n16343), .B2(n5675), .A(n5676), .ZN(n5673) );
  OAI21_X2 U8647 ( .B1(n16340), .B2(n5491), .A(n5492), .ZN(n5489) );
  OAI21_X2 U8648 ( .B1(n16326), .B2(n5312), .A(n5313), .ZN(n5310) );
  OAI21_X2 U8649 ( .B1(n16310), .B2(n5114), .A(n5115), .ZN(n5112) );
  OAI21_X2 U8650 ( .B1(n16307), .B2(n4864), .A(n4865), .ZN(n4862) );
  OAI21_X2 U8651 ( .B1(n16292), .B2(n4606), .A(n4607), .ZN(n4604) );
  OAI21_X2 U8652 ( .B1(n16280), .B2(n4325), .A(n4326), .ZN(n4323) );
  OAI21_X2 U8653 ( .B1(n16269), .B2(n4026), .A(n4027), .ZN(n4024) );
  OAI21_X2 U8654 ( .B1(n16265), .B2(n3722), .A(n3723), .ZN(n3720) );
  OAI21_X2 U8655 ( .B1(n16261), .B2(n3298), .A(n3299), .ZN(n3296) );
  OAI21_X2 U8656 ( .B1(n16259), .B2(n3290), .A(n3291), .ZN(n3288) );
  OAI21_X2 U8657 ( .B1(n5851), .B2(n5850), .A(n5871), .ZN(n5845) );
  OAI21_X2 U8658 ( .B1(n5764), .B2(n5765), .A(n5694), .ZN(n5763) );
  OAI21_X2 U8659 ( .B1(n5550), .B2(n5551), .A(n5525), .ZN(n5549) );
  OAI21_X2 U8660 ( .B1(n5178), .B2(n5179), .A(n5157), .ZN(n5177) );
  OAI21_X2 U8661 ( .B1(n5941), .B2(n5942), .A(n5943), .ZN(n5940) );
  OAI21_X2 U8662 ( .B1(n5863), .B2(n5864), .A(n5779), .ZN(n5862) );
  OAI21_X2 U8663 ( .B1(n5672), .B2(n5673), .A(n5607), .ZN(n5671) );
  OAI21_X2 U8664 ( .B1(n5488), .B2(n5489), .A(n5441), .ZN(n5487) );
  OAI21_X2 U8665 ( .B1(n5111), .B2(n5112), .A(n5050), .ZN(n5110) );
  OAI21_X2 U8666 ( .B1(n4861), .B2(n4862), .A(n4792), .ZN(n4860) );
  OAI21_X2 U8667 ( .B1(n4023), .B2(n4024), .A(n3941), .ZN(n4022) );
  OAI21_X2 U8668 ( .B1(n5231), .B2(n5232), .A(n5233), .ZN(n5230) );
  OAI21_X2 U8669 ( .B1(n16341), .B2(n5573), .A(n5574), .ZN(n5571) );
  OAI21_X2 U8670 ( .B1(n16328), .B2(n5484), .A(n5485), .ZN(n5482) );
  OAI21_X2 U8671 ( .B1(n5212), .B2(n5213), .A(n5214), .ZN(n5211) );
  OAI21_X2 U8672 ( .B1(n16309), .B2(n5107), .A(n5108), .ZN(n5105) );
  OAI21_X2 U8673 ( .B1(n16293), .B2(n4735), .A(n4736), .ZN(n4733) );
  OAI21_X2 U8674 ( .B1(n16303), .B2(n4851), .A(n4852), .ZN(n4849) );
  OAI21_X2 U8675 ( .B1(n16290), .B2(n4599), .A(n4600), .ZN(n4597) );
  OAI21_X2 U8676 ( .B1(n16297), .B2(n4839), .A(n4840), .ZN(n4837) );
  OAI21_X2 U8677 ( .B1(n16281), .B2(n4465), .A(n4466), .ZN(n4463) );
  OAI21_X2 U8678 ( .B1(n16287), .B2(n4717), .A(n4718), .ZN(n4715) );
  OAI21_X2 U8679 ( .B1(n16286), .B2(n4587), .A(n4588), .ZN(n4585) );
  OAI21_X2 U8680 ( .B1(n16270), .B2(n4173), .A(n4174), .ZN(n4171) );
  OAI21_X2 U8681 ( .B1(n5971), .B2(n5972), .A(n5973), .ZN(n5970) );
  OAI21_X2 U8682 ( .B1(n16302), .B2(n5190), .A(n5191), .ZN(n5188) );
  OAI21_X2 U8683 ( .B1(n16345), .B2(n5746), .A(n5747), .ZN(n5744) );
  OAI21_X2 U8684 ( .B1(n16327), .B2(n5402), .A(n5403), .ZN(n5400) );
  OAI21_X2 U8685 ( .B1(n3871), .B2(n3872), .A(n3873), .ZN(n3870) );
  OAI21_X2 U8686 ( .B1(n16342), .B2(n5668), .A(n5669), .ZN(n5666) );
  OAI21_X2 U8687 ( .B1(n5566), .B2(n5567), .A(n5568), .ZN(n5565) );
  OAI21_X2 U8688 ( .B1(n5477), .B2(n5478), .A(n5479), .ZN(n5476) );
  OAI21_X2 U8689 ( .B1(n5206), .B2(n5207), .A(n5208), .ZN(n5205) );
  OAI21_X2 U8690 ( .B1(n16301), .B2(n5089), .A(n5090), .ZN(n5087) );
  OAI21_X2 U8691 ( .B1(n4976), .B2(n4977), .A(n4978), .ZN(n4975) );
  OAI21_X2 U8692 ( .B1(n5751), .B2(n5752), .A(n5753), .ZN(n5750) );
  OAI21_X2 U8693 ( .B1(n16308), .B2(n5001), .A(n5002), .ZN(n4999) );
  OAI21_X2 U8694 ( .B1(n5100), .B2(n5101), .A(n5102), .ZN(n5099) );
  OAI21_X2 U8695 ( .B1(n16306), .B2(n4995), .A(n4996), .ZN(n4993) );
  OAI21_X2 U8696 ( .B1(n16305), .B2(n4857), .A(n4858), .ZN(n4855) );
  OAI21_X2 U8697 ( .B1(n16304), .B2(n4989), .A(n4990), .ZN(n4987) );
  OAI21_X2 U8698 ( .B1(n16300), .B2(n4983), .A(n4984), .ZN(n4981) );
  OAI21_X2 U8699 ( .B1(n16291), .B2(n4729), .A(n4730), .ZN(n4727) );
  OAI21_X2 U8700 ( .B1(n16299), .B2(n4845), .A(n4846), .ZN(n4843) );
  OAI21_X2 U8701 ( .B1(n16289), .B2(n4723), .A(n4724), .ZN(n4721) );
  OAI21_X2 U8702 ( .B1(n16288), .B2(n4593), .A(n4594), .ZN(n4591) );
  OAI21_X2 U8703 ( .B1(n16279), .B2(n4459), .A(n4460), .ZN(n4457) );
  OAI21_X2 U8704 ( .B1(n4832), .B2(n4833), .A(n4834), .ZN(n4831) );
  OAI21_X2 U8705 ( .B1(n16278), .B2(n4318), .A(n4319), .ZN(n4316) );
  OAI21_X2 U8706 ( .B1(n16285), .B2(n4711), .A(n4712), .ZN(n4709) );
  OAI21_X2 U8707 ( .B1(n16277), .B2(n4453), .A(n4454), .ZN(n4451) );
  OAI21_X2 U8708 ( .B1(n16284), .B2(n4581), .A(n4582), .ZN(n4579) );
  OAI21_X2 U8709 ( .B1(n16276), .B2(n4312), .A(n4313), .ZN(n4310) );
  OAI21_X2 U8710 ( .B1(n16275), .B2(n4447), .A(n4448), .ZN(n4445) );
  OAI21_X2 U8711 ( .B1(n16274), .B2(n4306), .A(n4307), .ZN(n4304) );
  OAI21_X2 U8712 ( .B1(n16339), .B2(n5346), .A(n5347), .ZN(n5344) );
  OAI21_X2 U8713 ( .B1(n5856), .B2(n5857), .A(n5858), .ZN(n5855) );
  OAI21_X2 U8714 ( .B1(n5820), .B2(n5821), .A(n5822), .ZN(n5819) );
  BUF_X4 U8715 ( .A(n12882), .Z(n13004) );
  BUF_X4 U8716 ( .A(n12898), .Z(n12954) );
  BUF_X4 U8717 ( .A(n12882), .Z(n13003) );
  BUF_X4 U8718 ( .A(n12882), .Z(n13002) );
  BUF_X4 U8719 ( .A(n12883), .Z(n13001) );
  BUF_X4 U8720 ( .A(n12883), .Z(n13000) );
  BUF_X4 U8721 ( .A(n12883), .Z(n12999) );
  BUF_X4 U8722 ( .A(n12899), .Z(n12953) );
  BUF_X4 U8723 ( .A(n12884), .Z(n12998) );
  BUF_X4 U8724 ( .A(n12900), .Z(n12948) );
  BUF_X4 U8725 ( .A(n12884), .Z(n12997) );
  BUF_X4 U8726 ( .A(n12884), .Z(n12996) );
  BUF_X4 U8727 ( .A(n12885), .Z(n12995) );
  BUF_X4 U8728 ( .A(n12885), .Z(n12994) );
  BUF_X4 U8729 ( .A(n12885), .Z(n12993) );
  BUF_X4 U8730 ( .A(n12901), .Z(n12947) );
  BUF_X4 U8731 ( .A(n12886), .Z(n12992) );
  BUF_X4 U8732 ( .A(n12886), .Z(n12991) );
  BUF_X4 U8733 ( .A(n13013), .Z(n13042) );
  BUF_X4 U8734 ( .A(n13006), .Z(n13060) );
  BUF_X4 U8735 ( .A(n13014), .Z(n13039) );
  BUF_X4 U8736 ( .A(n13007), .Z(n13059) );
  BUF_X4 U8737 ( .A(n13007), .Z(n13058) );
  BUF_X4 U8738 ( .A(n13007), .Z(n13057) );
  BUF_X4 U8739 ( .A(n12886), .Z(n12990) );
  BUF_X4 U8740 ( .A(n12902), .Z(n12944) );
  BUF_X4 U8741 ( .A(n12887), .Z(n12989) );
  BUF_X4 U8742 ( .A(n12902), .Z(n12943) );
  BUF_X4 U8743 ( .A(n12902), .Z(n12942) );
  BUF_X4 U8744 ( .A(n12887), .Z(n12988) );
  BUF_X4 U8745 ( .A(n12903), .Z(n12941) );
  BUF_X4 U8746 ( .A(n12889), .Z(n12983) );
  BUF_X4 U8747 ( .A(n12888), .Z(n12984) );
  BUF_X4 U8748 ( .A(n12904), .Z(n12938) );
  BUF_X4 U8749 ( .A(n12904), .Z(n12937) );
  BUF_X4 U8750 ( .A(n12887), .Z(n12987) );
  BUF_X4 U8751 ( .A(n12888), .Z(n12986) );
  BUF_X4 U8752 ( .A(n12888), .Z(n12985) );
  BUF_X4 U8753 ( .A(n12903), .Z(n12940) );
  BUF_X4 U8754 ( .A(n12903), .Z(n12939) );
  BUF_X4 U8755 ( .A(n12889), .Z(n12982) );
  BUF_X4 U8756 ( .A(n12904), .Z(n12936) );
  BUF_X4 U8757 ( .A(n12905), .Z(n12935) );
  BUF_X4 U8758 ( .A(n12891), .Z(n12977) );
  BUF_X4 U8759 ( .A(n12890), .Z(n12978) );
  BUF_X4 U8760 ( .A(n12906), .Z(n12932) );
  BUF_X4 U8761 ( .A(n12906), .Z(n12931) );
  BUF_X4 U8762 ( .A(n12889), .Z(n12981) );
  BUF_X4 U8763 ( .A(n12890), .Z(n12980) );
  BUF_X4 U8764 ( .A(n12890), .Z(n12979) );
  BUF_X4 U8765 ( .A(n12905), .Z(n12934) );
  BUF_X4 U8766 ( .A(n12905), .Z(n12933) );
  BUF_X4 U8767 ( .A(n12891), .Z(n12976) );
  BUF_X4 U8768 ( .A(n12906), .Z(n12930) );
  BUF_X4 U8769 ( .A(n12907), .Z(n12929) );
  BUF_X4 U8770 ( .A(n12908), .Z(n12925) );
  BUF_X4 U8771 ( .A(n12892), .Z(n12973) );
  BUF_X4 U8772 ( .A(n12892), .Z(n12972) );
  BUF_X4 U8773 ( .A(n12908), .Z(n12926) );
  BUF_X4 U8774 ( .A(n12891), .Z(n12975) );
  BUF_X4 U8775 ( .A(n12892), .Z(n12974) );
  BUF_X4 U8776 ( .A(n12907), .Z(n12928) );
  BUF_X4 U8777 ( .A(n12907), .Z(n12927) );
  BUF_X4 U8778 ( .A(n12912), .Z(n12913) );
  BUF_X4 U8779 ( .A(n12896), .Z(n12961) );
  BUF_X4 U8780 ( .A(n12896), .Z(n12960) );
  BUF_X4 U8781 ( .A(n12912), .Z(n12914) );
  BUF_X4 U8782 ( .A(n12895), .Z(n12964) );
  BUF_X4 U8783 ( .A(n12895), .Z(n12963) );
  BUF_X4 U8784 ( .A(n12896), .Z(n12962) );
  BUF_X4 U8785 ( .A(n12911), .Z(n12917) );
  BUF_X4 U8786 ( .A(n12911), .Z(n12916) );
  BUF_X4 U8787 ( .A(n12911), .Z(n12915) );
  BUF_X4 U8788 ( .A(n12895), .Z(n12965) );
  BUF_X4 U8789 ( .A(n12910), .Z(n12919) );
  BUF_X4 U8790 ( .A(n12910), .Z(n12918) );
  BUF_X4 U8791 ( .A(n12894), .Z(n12967) );
  BUF_X4 U8792 ( .A(n12894), .Z(n12966) );
  BUF_X4 U8793 ( .A(n12910), .Z(n12920) );
  BUF_X4 U8794 ( .A(n12893), .Z(n12971) );
  BUF_X4 U8795 ( .A(n12893), .Z(n12970) );
  BUF_X4 U8796 ( .A(n12908), .Z(n12924) );
  BUF_X4 U8797 ( .A(n12893), .Z(n12969) );
  BUF_X4 U8798 ( .A(n12894), .Z(n12968) );
  BUF_X4 U8799 ( .A(n12909), .Z(n12923) );
  BUF_X4 U8800 ( .A(n12909), .Z(n12922) );
  BUF_X4 U8801 ( .A(n12909), .Z(n12921) );
  BUF_X4 U8802 ( .A(n13015), .Z(n13036) );
  BUF_X4 U8803 ( .A(n13008), .Z(n13056) );
  BUF_X4 U8804 ( .A(n13008), .Z(n13055) );
  BUF_X4 U8805 ( .A(n13016), .Z(n13035) );
  BUF_X4 U8806 ( .A(n13016), .Z(n13034) );
  BUF_X4 U8807 ( .A(n13009), .Z(n13054) );
  BUF_X4 U8808 ( .A(n13016), .Z(n13033) );
  BUF_X4 U8809 ( .A(n13009), .Z(n13053) );
  BUF_X4 U8810 ( .A(n13009), .Z(n13052) );
  BUF_X4 U8811 ( .A(n13017), .Z(n13032) );
  BUF_X4 U8812 ( .A(n13017), .Z(n13031) );
  BUF_X4 U8813 ( .A(n13017), .Z(n13030) );
  BUF_X4 U8814 ( .A(n13010), .Z(n13050) );
  BUF_X4 U8815 ( .A(n13010), .Z(n13051) );
  BUF_X4 U8816 ( .A(n13018), .Z(n13029) );
  BUF_X4 U8817 ( .A(n13018), .Z(n13028) );
  BUF_X4 U8818 ( .A(n13012), .Z(n13044) );
  BUF_X4 U8819 ( .A(n13012), .Z(n13045) );
  BUF_X4 U8820 ( .A(n13020), .Z(n13023) );
  BUF_X4 U8821 ( .A(n13020), .Z(n13022) );
  BUF_X4 U8822 ( .A(n13012), .Z(n13046) );
  BUF_X4 U8823 ( .A(n13019), .Z(n13024) );
  BUF_X4 U8824 ( .A(n13011), .Z(n13047) );
  BUF_X4 U8825 ( .A(n13011), .Z(n13049) );
  BUF_X4 U8826 ( .A(n13018), .Z(n13027) );
  BUF_X4 U8827 ( .A(n13011), .Z(n13048) );
  BUF_X4 U8828 ( .A(n13019), .Z(n13026) );
  BUF_X4 U8829 ( .A(n13019), .Z(n13025) );
  BUF_X4 U8830 ( .A(n12897), .Z(n12959) );
  BUF_X4 U8831 ( .A(n12897), .Z(n12958) );
  BUF_X4 U8832 ( .A(n12897), .Z(n12957) );
  BUF_X4 U8833 ( .A(n12898), .Z(n12956) );
  BUF_X4 U8834 ( .A(n12898), .Z(n12955) );
  BUF_X4 U8835 ( .A(n12899), .Z(n12952) );
  BUF_X4 U8836 ( .A(n12899), .Z(n12951) );
  BUF_X4 U8837 ( .A(n12900), .Z(n12950) );
  BUF_X4 U8838 ( .A(n12900), .Z(n12949) );
  BUF_X4 U8839 ( .A(n12901), .Z(n12946) );
  BUF_X4 U8840 ( .A(n12901), .Z(n12945) );
  BUF_X4 U8841 ( .A(n13013), .Z(n13043) );
  BUF_X4 U8842 ( .A(n13014), .Z(n13041) );
  BUF_X4 U8843 ( .A(n13014), .Z(n13040) );
  BUF_X4 U8844 ( .A(n13015), .Z(n13038) );
  BUF_X4 U8845 ( .A(n13015), .Z(n13037) );
  BUF_X4 U8846 ( .A(n10757), .Z(n10834) );
  BUF_X4 U8847 ( .A(n10757), .Z(n10833) );
  BUF_X4 U8848 ( .A(n10773), .Z(n10787) );
  BUF_X4 U8849 ( .A(n10773), .Z(n10786) );
  BUF_X4 U8850 ( .A(n10775), .Z(n10780) );
  BUF_X4 U8851 ( .A(n10760), .Z(n10826) );
  BUF_X4 U8852 ( .A(n10760), .Z(n10825) );
  BUF_X4 U8853 ( .A(n10775), .Z(n10779) );
  BUF_X4 U8854 ( .A(n10761), .Z(n10821) );
  BUF_X4 U8855 ( .A(n10752), .Z(n10850) );
  BUF_X4 U8856 ( .A(n10757), .Z(n10835) );
  BUF_X4 U8857 ( .A(n10772), .Z(n10789) );
  BUF_X4 U8858 ( .A(n10772), .Z(n10788) );
  BUF_X4 U8859 ( .A(n10762), .Z(n10820) );
  BUF_X4 U8860 ( .A(n10748), .Z(n10861) );
  BUF_X4 U8861 ( .A(n10763), .Z(n10816) );
  BUF_X4 U8862 ( .A(n10763), .Z(n10815) );
  BUF_X4 U8863 ( .A(n10748), .Z(n10860) );
  BUF_X4 U8864 ( .A(n10748), .Z(n10859) );
  BUF_X4 U8865 ( .A(n10764), .Z(n10814) );
  BUF_X4 U8866 ( .A(n10751), .Z(n10853) );
  BUF_X4 U8867 ( .A(n10766), .Z(n10806) );
  BUF_X4 U8868 ( .A(n10764), .Z(n10813) );
  BUF_X4 U8869 ( .A(n10764), .Z(n10812) );
  BUF_X4 U8870 ( .A(n10749), .Z(n10858) );
  BUF_X4 U8871 ( .A(n10749), .Z(n10857) );
  BUF_X4 U8872 ( .A(n10765), .Z(n10811) );
  BUF_X4 U8873 ( .A(n10750), .Z(n10856) );
  BUF_X4 U8874 ( .A(n10765), .Z(n10810) );
  BUF_X4 U8875 ( .A(n10765), .Z(n10809) );
  BUF_X4 U8876 ( .A(n10750), .Z(n10855) );
  BUF_X4 U8877 ( .A(n10750), .Z(n10854) );
  BUF_X4 U8878 ( .A(n10766), .Z(n10808) );
  BUF_X4 U8879 ( .A(n10766), .Z(n10807) );
  BUF_X4 U8880 ( .A(n10769), .Z(n10799) );
  BUF_X4 U8881 ( .A(n10756), .Z(n10837) );
  BUF_X4 U8882 ( .A(n10756), .Z(n10836) );
  BUF_X4 U8883 ( .A(n10772), .Z(n10790) );
  BUF_X4 U8884 ( .A(n10758), .Z(n10832) );
  BUF_X4 U8885 ( .A(n10758), .Z(n10831) );
  BUF_X4 U8886 ( .A(n10773), .Z(n10785) );
  BUF_X4 U8887 ( .A(n10770), .Z(n10796) );
  BUF_X4 U8888 ( .A(n10771), .Z(n10793) );
  BUF_X4 U8889 ( .A(n10758), .Z(n10830) );
  BUF_X4 U8890 ( .A(n10774), .Z(n10784) );
  BUF_X4 U8891 ( .A(n10774), .Z(n10783) );
  BUF_X4 U8892 ( .A(n10759), .Z(n10829) );
  BUF_X4 U8893 ( .A(n10759), .Z(n10828) );
  BUF_X4 U8894 ( .A(n10759), .Z(n10827) );
  BUF_X4 U8895 ( .A(n10774), .Z(n10782) );
  BUF_X4 U8896 ( .A(n10775), .Z(n10781) );
  BUF_X4 U8897 ( .A(n10753), .Z(n10847) );
  BUF_X4 U8898 ( .A(n10753), .Z(n10846) );
  BUF_X4 U8899 ( .A(n10768), .Z(n10800) );
  BUF_X4 U8900 ( .A(n10753), .Z(n10845) );
  BUF_X4 U8901 ( .A(n10754), .Z(n10844) );
  BUF_X4 U8902 ( .A(n10754), .Z(n10843) );
  BUF_X4 U8903 ( .A(n10769), .Z(n10798) );
  BUF_X4 U8904 ( .A(n10769), .Z(n10797) );
  BUF_X4 U8905 ( .A(n10754), .Z(n10842) );
  BUF_X4 U8906 ( .A(n10755), .Z(n10841) );
  BUF_X4 U8907 ( .A(n10755), .Z(n10840) );
  BUF_X4 U8908 ( .A(n10770), .Z(n10795) );
  BUF_X4 U8909 ( .A(n10770), .Z(n10794) );
  BUF_X4 U8910 ( .A(n10755), .Z(n10839) );
  BUF_X4 U8911 ( .A(n10756), .Z(n10838) );
  BUF_X4 U8912 ( .A(n10771), .Z(n10792) );
  BUF_X4 U8913 ( .A(n10771), .Z(n10791) );
  BUF_X4 U8914 ( .A(n10747), .Z(n10862) );
  BUF_X4 U8915 ( .A(n10762), .Z(n10819) );
  BUF_X4 U8916 ( .A(n10762), .Z(n10818) );
  BUF_X4 U8917 ( .A(n10763), .Z(n10817) );
  BUF_X4 U8918 ( .A(n10760), .Z(n10824) );
  BUF_X4 U8919 ( .A(n10776), .Z(n10778) );
  BUF_X4 U8920 ( .A(n10776), .Z(n10777) );
  BUF_X4 U8921 ( .A(n10761), .Z(n10823) );
  BUF_X4 U8922 ( .A(n10761), .Z(n10822) );
  BUF_X4 U8923 ( .A(n10751), .Z(n10852) );
  BUF_X4 U8924 ( .A(n10751), .Z(n10851) );
  BUF_X4 U8925 ( .A(n10767), .Z(n10805) );
  BUF_X4 U8926 ( .A(n10767), .Z(n10804) );
  BUF_X4 U8927 ( .A(n10752), .Z(n10849) );
  BUF_X4 U8928 ( .A(n10752), .Z(n10848) );
  BUF_X4 U8929 ( .A(n10767), .Z(n10803) );
  BUF_X4 U8930 ( .A(n10768), .Z(n10802) );
  BUF_X4 U8931 ( .A(n10768), .Z(n10801) );
  BUF_X4 U8932 ( .A(n13020), .Z(n13021) );
  INV_X4 U8933 ( .A(n13096), .ZN(n13101) );
  INV_X4 U8934 ( .A(n13096), .ZN(n13098) );
  INV_X4 U8935 ( .A(n13096), .ZN(n13100) );
  INV_X4 U8936 ( .A(n13096), .ZN(n13097) );
  INV_X4 U8937 ( .A(n13096), .ZN(n13099) );
  INV_X4 U8938 ( .A(n13095), .ZN(n13092) );
  INV_X4 U8939 ( .A(n13095), .ZN(n13094) );
  INV_X4 U8940 ( .A(n13095), .ZN(n13093) );
  NAND2_X2 U8941 ( .A1(n16456), .A2(n16469), .ZN(n3964) );
  BUF_X4 U8942 ( .A(n10877), .Z(n10884) );
  BUF_X4 U8943 ( .A(n10869), .Z(n10908) );
  BUF_X4 U8944 ( .A(n10876), .Z(n10885) );
  BUF_X4 U8945 ( .A(n10871), .Z(n10901) );
  BUF_X4 U8946 ( .A(n10864), .Z(n10920) );
  BUF_X4 U8947 ( .A(n10872), .Z(n10898) );
  BUF_X4 U8948 ( .A(n10872), .Z(n10897) );
  BUF_X4 U8949 ( .A(n10865), .Z(n10919) );
  BUF_X4 U8950 ( .A(n10873), .Z(n10896) );
  BUF_X4 U8951 ( .A(n10865), .Z(n10918) );
  BUF_X4 U8952 ( .A(n10873), .Z(n10895) );
  BUF_X4 U8953 ( .A(n10873), .Z(n10894) );
  BUF_X4 U8954 ( .A(n10868), .Z(n10909) );
  BUF_X4 U8955 ( .A(n10869), .Z(n10907) );
  BUF_X4 U8956 ( .A(n10869), .Z(n10906) );
  BUF_X4 U8957 ( .A(n10877), .Z(n10883) );
  BUF_X4 U8958 ( .A(n10870), .Z(n10905) );
  BUF_X4 U8959 ( .A(n10870), .Z(n10904) );
  BUF_X4 U8960 ( .A(n10877), .Z(n10882) );
  BUF_X4 U8961 ( .A(n10878), .Z(n10881) );
  BUF_X4 U8962 ( .A(n10867), .Z(n10914) );
  BUF_X4 U8963 ( .A(n10867), .Z(n10913) );
  BUF_X4 U8964 ( .A(n10875), .Z(n10890) );
  BUF_X4 U8965 ( .A(n10875), .Z(n10889) );
  BUF_X4 U8966 ( .A(n10867), .Z(n10912) );
  BUF_X4 U8967 ( .A(n10868), .Z(n10911) );
  BUF_X4 U8968 ( .A(n10875), .Z(n10888) );
  BUF_X4 U8969 ( .A(n10868), .Z(n10910) );
  BUF_X4 U8970 ( .A(n10876), .Z(n10887) );
  BUF_X4 U8971 ( .A(n10876), .Z(n10886) );
  BUF_X4 U8972 ( .A(n10871), .Z(n10900) );
  BUF_X4 U8973 ( .A(n10872), .Z(n10899) );
  BUF_X4 U8974 ( .A(n10870), .Z(n10903) );
  BUF_X4 U8975 ( .A(n10878), .Z(n10880) );
  BUF_X4 U8976 ( .A(n10871), .Z(n10902) );
  BUF_X4 U8977 ( .A(n10866), .Z(n10917) );
  BUF_X4 U8978 ( .A(n10866), .Z(n10916) );
  BUF_X4 U8979 ( .A(n10874), .Z(n10893) );
  BUF_X4 U8980 ( .A(n10866), .Z(n10915) );
  BUF_X4 U8981 ( .A(n10874), .Z(n10892) );
  BUF_X4 U8982 ( .A(n10874), .Z(n10891) );
  BUF_X4 U8983 ( .A(n10878), .Z(n10879) );
  INV_X4 U8984 ( .A(n8807), .ZN(n13226) );
  INV_X4 U8985 ( .A(n8808), .ZN(n13106) );
  INV_X4 U8986 ( .A(n8808), .ZN(n13105) );
  INV_X4 U8987 ( .A(decode_rs2_4_), .ZN(n10955) );
  INV_X4 U8988 ( .A(n8807), .ZN(n13227) );
  INV_X4 U8989 ( .A(n13223), .ZN(n13222) );
  INV_X4 U8990 ( .A(n13223), .ZN(n13221) );
  INV_X4 U8991 ( .A(n8662), .ZN(n13506) );
  INV_X4 U8992 ( .A(n8662), .ZN(n13505) );
  INV_X4 U8993 ( .A(n8698), .ZN(n13511) );
  INV_X4 U8994 ( .A(n8698), .ZN(n13510) );
  INV_X4 U8995 ( .A(n8663), .ZN(n13516) );
  INV_X4 U8996 ( .A(n8663), .ZN(n13515) );
  INV_X4 U8997 ( .A(n8664), .ZN(n13521) );
  INV_X4 U8998 ( .A(n8664), .ZN(n13520) );
  INV_X4 U8999 ( .A(n8662), .ZN(n13507) );
  INV_X4 U9000 ( .A(n8698), .ZN(n13512) );
  INV_X4 U9001 ( .A(n8663), .ZN(n13517) );
  INV_X4 U9002 ( .A(n8664), .ZN(n13522) );
  INV_X4 U9003 ( .A(n8662), .ZN(n13508) );
  INV_X4 U9004 ( .A(n8698), .ZN(n13513) );
  INV_X4 U9005 ( .A(n8663), .ZN(n13518) );
  INV_X4 U9006 ( .A(n8664), .ZN(n13523) );
  INV_X4 U9007 ( .A(n8662), .ZN(n13509) );
  INV_X4 U9008 ( .A(n8698), .ZN(n13514) );
  INV_X4 U9009 ( .A(n8663), .ZN(n13519) );
  INV_X4 U9010 ( .A(n8664), .ZN(n13524) );
  AOI21_X2 U9011 ( .B1(n5661), .B2(n5662), .A(n5663), .ZN(n5566) );
  AOI21_X2 U9012 ( .B1(n5560), .B2(n5561), .A(n5562), .ZN(n5477) );
  AOI21_X2 U9013 ( .B1(n5471), .B2(n5472), .A(n5473), .ZN(n5390) );
  AOI21_X2 U9014 ( .B1(n5299), .B2(n5300), .A(n5301), .ZN(n5206) );
  AOI21_X2 U9015 ( .B1(n5082), .B2(n5083), .A(n5084), .ZN(n4976) );
  AOI21_X2 U9016 ( .B1(n3988), .B2(n3989), .A(n3990), .ZN(n3840) );
  AOI21_X2 U9017 ( .B1(n3689), .B2(n3690), .A(n3691), .ZN(n3503) );
  AOI21_X2 U9018 ( .B1(n5912), .B2(n5913), .A(n5914), .ZN(n5894) );
  AOI21_X2 U9019 ( .B1(n5877), .B2(n5878), .A(n16348), .ZN(n5851) );
  AOI21_X2 U9020 ( .B1(n5304), .B2(n5305), .A(n5306), .ZN(n5212) );
  AOI21_X2 U9021 ( .B1(n5385), .B2(n5386), .A(n5387), .ZN(n5294) );
  AOI21_X2 U9022 ( .B1(n5380), .B2(n5381), .A(n5382), .ZN(n5289) );
  AOI21_X2 U9023 ( .B1(n5200), .B2(n5201), .A(n5202), .ZN(n5100) );
  AOI21_X2 U9024 ( .B1(n4970), .B2(n4971), .A(n4972), .ZN(n4832) );
  AOI21_X2 U9025 ( .B1(n4028), .B2(n4029), .A(n4030), .ZN(n3878) );
  AOI21_X2 U9026 ( .B1(n4698), .B2(n4699), .A(n4700), .ZN(n4568) );
  AOI21_X2 U9027 ( .B1(n4018), .B2(n4019), .A(n4020), .ZN(n3871) );
  AOI21_X2 U9028 ( .B1(n4013), .B2(n4014), .A(n4015), .ZN(n3865) );
  AOI21_X2 U9029 ( .B1(n4008), .B2(n4009), .A(n4010), .ZN(n3860) );
  AOI21_X2 U9030 ( .B1(n3709), .B2(n3710), .A(n3711), .ZN(n3532) );
  AOI21_X2 U9031 ( .B1(n3998), .B2(n3999), .A(n4000), .ZN(n3850) );
  AOI21_X2 U9032 ( .B1(n3704), .B2(n3705), .A(n3706), .ZN(n3524) );
  AOI21_X2 U9033 ( .B1(n3993), .B2(n3994), .A(n3995), .ZN(n3845) );
  AOI21_X2 U9034 ( .B1(n3699), .B2(n3700), .A(n3701), .ZN(n3518) );
  AOI21_X2 U9035 ( .B1(n4131), .B2(n4132), .A(n4133), .ZN(n3983) );
  AOI21_X2 U9036 ( .B1(n3835), .B2(n3836), .A(n3837), .ZN(n3684) );
  AOI21_X2 U9037 ( .B1(n4126), .B2(n4127), .A(n4128), .ZN(n3978) );
  AOI21_X2 U9038 ( .B1(n3496), .B2(n3497), .A(n3498), .ZN(n3271) );
  AOI21_X2 U9039 ( .B1(n3489), .B2(n3490), .A(n3491), .ZN(n3375) );
  AOI21_X2 U9040 ( .B1(n3462), .B2(n3463), .A(n3464), .ZN(n3382) );
  AOI21_X2 U9041 ( .B1(n5282), .B2(n5283), .A(n5284), .ZN(n5183) );
  AOI21_X2 U9042 ( .B1(n5884), .B2(n5883), .A(n5931), .ZN(n5887) );
  AOI21_X2 U9043 ( .B1(n5904), .B2(n5905), .A(n5906), .ZN(n5771) );
  AOI21_X2 U9044 ( .B1(n5869), .B2(n5870), .A(n5907), .ZN(n5774) );
  AOI21_X2 U9045 ( .B1(n5511), .B2(n5512), .A(n5513), .ZN(n5427) );
  AOI21_X2 U9046 ( .B1(n5698), .B2(n5699), .A(n5700), .ZN(n5599) );
  AOI21_X2 U9047 ( .B1(n5514), .B2(n5515), .A(n5516), .ZN(n5430) );
  AOI21_X2 U9048 ( .B1(n5701), .B2(n5702), .A(n5703), .ZN(n5602) );
  AOI21_X2 U9049 ( .B1(n5335), .B2(n5336), .A(n5337), .ZN(n5246) );
  AOI21_X2 U9050 ( .B1(n5520), .B2(n5521), .A(n5522), .ZN(n5436) );
  AOI21_X2 U9051 ( .B1(n5338), .B2(n5339), .A(n5340), .ZN(n5249) );
  AOI21_X2 U9052 ( .B1(n5140), .B2(n5141), .A(n5142), .ZN(n5033) );
  AOI21_X2 U9053 ( .B1(n5341), .B2(n5342), .A(n5343), .ZN(n5252) );
  AOI21_X2 U9054 ( .B1(n5146), .B2(n5147), .A(n5148), .ZN(n5039) );
  AOI21_X2 U9055 ( .B1(n5149), .B2(n5150), .A(n5151), .ZN(n5042) );
  AOI21_X2 U9056 ( .B1(n4899), .B2(n4900), .A(n4901), .ZN(n4778) );
  AOI21_X2 U9057 ( .B1(n5152), .B2(n5153), .A(n5154), .ZN(n5045) );
  AOI21_X2 U9058 ( .B1(n4905), .B2(n4906), .A(n4907), .ZN(n4784) );
  AOI21_X2 U9059 ( .B1(n4908), .B2(n4909), .A(n4910), .ZN(n4787) );
  AOI21_X2 U9060 ( .B1(n4652), .B2(n4653), .A(n4654), .ZN(n4513) );
  AOI21_X2 U9061 ( .B1(n4658), .B2(n4659), .A(n4660), .ZN(n4519) );
  AOI21_X2 U9062 ( .B1(n4380), .B2(n4381), .A(n4382), .ZN(n4231) );
  AOI21_X2 U9063 ( .B1(n5508), .B2(n5509), .A(n5510), .ZN(n5424) );
  AOI21_X2 U9064 ( .B1(n5329), .B2(n5330), .A(n5331), .ZN(n5231) );
  NOR2_X2 U9065 ( .A1(n2963), .A2(n2964), .ZN(n2962) );
  OAI21_X2 U9066 ( .B1(n5977), .B2(n5978), .A(n5979), .ZN(n5975) );
  OAI21_X2 U9067 ( .B1(n6001), .B2(n6002), .A(n5921), .ZN(n5999) );
  NOR3_X2 U9068 ( .A1(n2804), .A2(n13789), .A3(n5844), .ZN(n5841) );
  NOR3_X2 U9069 ( .A1(n13138), .A2(n2869), .A3(n5229), .ZN(n5139) );
  NOR3_X2 U9070 ( .A1(n13141), .A2(n13172), .A3(n5587), .ZN(n5510) );
  NOR3_X2 U9071 ( .A1(n8710), .A2(n13172), .A3(n5418), .ZN(n5331) );
  NOR3_X2 U9072 ( .A1(n13140), .A2(n13172), .A3(n5975), .ZN(n5974) );
  NOR3_X2 U9073 ( .A1(n13153), .A2(n13172), .A3(n5999), .ZN(n5914) );
  OAI21_X2 U9074 ( .B1(n13150), .B2(n13201), .A(n5956), .ZN(n5955) );
  OAI21_X2 U9075 ( .B1(n2775), .B2(n13148), .A(n5407), .ZN(n5406) );
  OAI21_X2 U9076 ( .B1(n13789), .B2(n3548), .A(n5288), .ZN(n5287) );
  OAI21_X2 U9077 ( .B1(n13159), .B2(n13139), .A(n4040), .ZN(n4039) );
  OAI21_X2 U9078 ( .B1(n3548), .B2(n13139), .A(n3549), .ZN(n3547) );
  OAI21_X2 U9079 ( .B1(n2869), .B2(n13155), .A(n5892), .ZN(n5891) );
  OAI21_X2 U9080 ( .B1(n2869), .B2(n13141), .A(n5500), .ZN(n5499) );
  OAI21_X2 U9081 ( .B1(n13189), .B2(n13148), .A(n5680), .ZN(n5679) );
  OAI21_X2 U9082 ( .B1(n13173), .B2(n13138), .A(n5325), .ZN(n5324) );
  OAI21_X2 U9083 ( .B1(n2830), .B2(n13146), .A(n5496), .ZN(n5495) );
  OAI21_X2 U9084 ( .B1(n2909), .B2(n13137), .A(n5321), .ZN(n5320) );
  OAI21_X2 U9085 ( .B1(n2804), .B2(n13148), .A(n5494), .ZN(n5493) );
  OAI21_X2 U9086 ( .B1(n2830), .B2(n13141), .A(n5319), .ZN(n5318) );
  OAI21_X2 U9087 ( .B1(n2804), .B2(n13135), .A(n5317), .ZN(n5316) );
  OAI21_X2 U9088 ( .B1(n2830), .B2(n8710), .A(n5123), .ZN(n5122) );
  OAI21_X2 U9089 ( .B1(n2909), .B2(n13139), .A(n4877), .ZN(n4876) );
  OAI21_X2 U9090 ( .B1(n2775), .B2(n13146), .A(n5315), .ZN(n5314) );
  OAI21_X2 U9091 ( .B1(n2804), .B2(n13137), .A(n5121), .ZN(n5120) );
  OAI21_X2 U9092 ( .B1(n2775), .B2(n13141), .A(n5119), .ZN(n5118) );
  OAI21_X2 U9093 ( .B1(n2804), .B2(n13138), .A(n4873), .ZN(n4872) );
  OAI21_X2 U9094 ( .B1(n2748), .B2(n13135), .A(n5117), .ZN(n5116) );
  OAI21_X2 U9095 ( .B1(n2804), .B2(n13139), .A(n4618), .ZN(n4617) );
  OAI21_X2 U9096 ( .B1(n2748), .B2(n13137), .A(n4869), .ZN(n4868) );
  OAI21_X2 U9097 ( .B1(n3569), .B2(n13141), .A(n4867), .ZN(n4866) );
  OAI21_X2 U9098 ( .B1(n2748), .B2(n13138), .A(n4614), .ZN(n4613) );
  OAI21_X2 U9099 ( .B1(n3569), .B2(n8710), .A(n4612), .ZN(n4611) );
  OAI21_X2 U9100 ( .B1(n2748), .B2(n13139), .A(n4337), .ZN(n4336) );
  OAI21_X2 U9101 ( .B1(n3565), .B2(n13137), .A(n4610), .ZN(n4609) );
  OAI21_X2 U9102 ( .B1(n3565), .B2(n13138), .A(n4333), .ZN(n4332) );
  OAI21_X2 U9103 ( .B1(n13180), .B2(n13138), .A(n4180), .ZN(n4179) );
  OAI21_X2 U9104 ( .B1(n13173), .B2(n13146), .A(n5763), .ZN(n5762) );
  OAI21_X2 U9105 ( .B1(n13172), .B2(n13137), .A(n5502), .ZN(n5501) );
  OAI21_X2 U9106 ( .B1(n13140), .B2(n2748), .A(n5665), .ZN(n5664) );
  OAI21_X2 U9107 ( .B1(n8738), .B2(n3569), .A(n5564), .ZN(n5563) );
  OAI21_X2 U9108 ( .B1(n13150), .B2(n13180), .A(n5653), .ZN(n5652) );
  OAI21_X2 U9109 ( .B1(n8738), .B2(n3565), .A(n5475), .ZN(n5474) );
  OAI21_X2 U9110 ( .B1(n13153), .B2(n3565), .A(n5303), .ZN(n5302) );
  OAI21_X2 U9111 ( .B1(n8738), .B2(n3548), .A(n5194), .ZN(n5193) );
  OAI21_X2 U9112 ( .B1(n13150), .B2(n13167), .A(n5281), .ZN(n5280) );
  OAI21_X2 U9113 ( .B1(n13140), .B2(n3293), .A(n5086), .ZN(n5085) );
  OAI21_X2 U9114 ( .B1(n13180), .B2(n13139), .A(n3887), .ZN(n3886) );
  OAI21_X2 U9115 ( .B1(n13137), .B2(n3548), .A(n4176), .ZN(n4175) );
  OAI21_X2 U9116 ( .B1(n8710), .B2(n3293), .A(n3875), .ZN(n3874) );
  OAI21_X2 U9117 ( .B1(n13138), .B2(n13167), .A(n3544), .ZN(n3541) );
  OAI21_X2 U9118 ( .B1(n2869), .B2(n13143), .A(n5966), .ZN(n5965) );
  OAI21_X2 U9119 ( .B1(n13142), .B2(n13209), .A(n5755), .ZN(n5754) );
  OAI21_X2 U9120 ( .B1(n13789), .B2(n2775), .A(n5840), .ZN(n5839) );
  OAI21_X2 U9121 ( .B1(n13153), .B2(n13212), .A(n5576), .ZN(n5575) );
  OAI21_X2 U9122 ( .B1(n13142), .B2(n2748), .A(n5570), .ZN(n5569) );
  OAI21_X2 U9123 ( .B1(n13142), .B2(n13157), .A(n5481), .ZN(n5480) );
  OAI21_X2 U9124 ( .B1(n13147), .B2(n3569), .A(n5216), .ZN(n5215) );
  OAI21_X2 U9125 ( .B1(n8738), .B2(n13180), .A(n5389), .ZN(n5388) );
  OAI21_X2 U9126 ( .B1(n8739), .B2(n3565), .A(n5210), .ZN(n5209) );
  OAI21_X2 U9127 ( .B1(n13151), .B2(n3548), .A(n5463), .ZN(n5462) );
  OAI21_X2 U9128 ( .B1(n13153), .B2(n13180), .A(n5204), .ZN(n5203) );
  OAI21_X2 U9129 ( .B1(n13145), .B2(n13159), .A(n5004), .ZN(n5003) );
  OAI21_X2 U9130 ( .B1(n8739), .B2(n13180), .A(n5104), .ZN(n5103) );
  OAI21_X2 U9131 ( .B1(n13142), .B2(n3555), .A(n5199), .ZN(n5198) );
  OAI21_X2 U9132 ( .B1(n13147), .B2(n13180), .A(n4998), .ZN(n4997) );
  OAI21_X2 U9133 ( .B1(n13154), .B2(n3555), .A(n5098), .ZN(n5097) );
  OAI21_X2 U9134 ( .B1(n8739), .B2(n3555), .A(n4992), .ZN(n4991) );
  OAI21_X2 U9135 ( .B1(n13142), .B2(n3548), .A(n5092), .ZN(n5091) );
  OAI21_X2 U9136 ( .B1(n13135), .B2(n13180), .A(n4738), .ZN(n4737) );
  OAI21_X2 U9137 ( .B1(n13147), .B2(n3555), .A(n4854), .ZN(n4853) );
  OAI21_X2 U9138 ( .B1(n13154), .B2(n3548), .A(n4986), .ZN(n4985) );
  OAI21_X2 U9139 ( .B1(n13145), .B2(n3555), .A(n4732), .ZN(n4731) );
  OAI21_X2 U9140 ( .B1(n8739), .B2(n13165), .A(n4848), .ZN(n4847) );
  OAI21_X2 U9141 ( .B1(n13142), .B2(n3293), .A(n4980), .ZN(n4979) );
  OAI21_X2 U9142 ( .B1(n13147), .B2(n3548), .A(n4726), .ZN(n4725) );
  OAI21_X2 U9143 ( .B1(n13180), .B2(n8710), .A(n4331), .ZN(n4330) );
  OAI21_X2 U9144 ( .B1(n13154), .B2(n3293), .A(n4842), .ZN(n4841) );
  OAI21_X2 U9145 ( .B1(n13141), .B2(n3555), .A(n4468), .ZN(n4467) );
  OAI21_X2 U9146 ( .B1(n13145), .B2(n3548), .A(n4596), .ZN(n4595) );
  OAI21_X2 U9147 ( .B1(n13140), .B2(n13167), .A(n4974), .ZN(n4973) );
  OAI21_X2 U9148 ( .B1(n8739), .B2(n3293), .A(n4720), .ZN(n4719) );
  OAI21_X2 U9149 ( .B1(n13135), .B2(n3548), .A(n4462), .ZN(n4461) );
  OAI21_X2 U9150 ( .B1(n13142), .B2(n13167), .A(n4836), .ZN(n4835) );
  OAI21_X2 U9151 ( .B1(n13147), .B2(n3293), .A(n4590), .ZN(n4589) );
  OAI21_X2 U9152 ( .B1(n13153), .B2(n13167), .A(n4714), .ZN(n4713) );
  OAI21_X2 U9153 ( .B1(n3555), .B2(n13138), .A(n4032), .ZN(n4031) );
  OAI21_X2 U9154 ( .B1(n13145), .B2(n13178), .A(n4456), .ZN(n4455) );
  OAI21_X2 U9155 ( .B1(n8739), .B2(n13167), .A(n4584), .ZN(n4583) );
  OAI21_X2 U9156 ( .B1(n13135), .B2(n3293), .A(n4315), .ZN(n4314) );
  OAI21_X2 U9157 ( .B1(n13147), .B2(n13167), .A(n4450), .ZN(n4449) );
  OAI21_X2 U9158 ( .B1(n13162), .B2(n13139), .A(n3733), .ZN(n3732) );
  OAI21_X2 U9159 ( .B1(n13145), .B2(n13167), .A(n4309), .ZN(n4308) );
  OAI21_X2 U9160 ( .B1(n13141), .B2(n13167), .A(n4017), .ZN(n4016) );
  OAI21_X2 U9161 ( .B1(n13172), .B2(n13135), .A(n5689), .ZN(n5688) );
  OAI21_X2 U9162 ( .B1(n13142), .B2(n2775), .A(n5671), .ZN(n5670) );
  OAI21_X2 U9163 ( .B1(n8739), .B2(n3569), .A(n5308), .ZN(n5307) );
  OAI21_X2 U9164 ( .B1(n13151), .B2(n3555), .A(n5549), .ZN(n5548) );
  OAI21_X2 U9165 ( .B1(n13147), .B2(n3565), .A(n5110), .ZN(n5109) );
  OAI21_X2 U9166 ( .B1(n13145), .B2(n13180), .A(n4860), .ZN(n4859) );
  OAI21_X2 U9167 ( .B1(n13135), .B2(n3555), .A(n4602), .ZN(n4601) );
  OAI21_X2 U9168 ( .B1(n13141), .B2(n3548), .A(n4321), .ZN(n4320) );
  OAI21_X2 U9169 ( .B1(n13137), .B2(n13178), .A(n4022), .ZN(n4021) );
  OAI21_X2 U9170 ( .B1(n8710), .B2(n13167), .A(n3718), .ZN(n3717) );
  OAI21_X2 U9171 ( .B1(n5588), .B2(n5589), .A(n5507), .ZN(n5587) );
  OAI21_X2 U9172 ( .B1(n5419), .B2(n5420), .A(n5328), .ZN(n5418) );
  OAI21_X2 U9173 ( .B1(n5962), .B2(n5961), .A(n5980), .ZN(n5964) );
  OAI21_X2 U9174 ( .B1(n4818), .B2(n4819), .A(n4820), .ZN(n4693) );
  OAI21_X2 U9175 ( .B1(n5075), .B2(n5076), .A(n5077), .ZN(n4965) );
  OAI21_X2 U9176 ( .B1(n5464), .B2(n5465), .A(n5466), .ZN(n5380) );
  OAI21_X2 U9177 ( .B1(n16266), .B2(n4157), .A(n4158), .ZN(n4008) );
  OAI21_X2 U9178 ( .B1(n3860), .B2(n3861), .A(n3862), .ZN(n3709) );
  OAI21_X2 U9179 ( .B1(n16203), .B2(n4147), .A(n4148), .ZN(n3998) );
  OAI21_X2 U9180 ( .B1(n3850), .B2(n3851), .A(n3852), .ZN(n3699) );
  OAI21_X2 U9181 ( .B1(n5739), .B2(n5740), .A(n5741), .ZN(n5661) );
  OAI21_X2 U9182 ( .B1(n5555), .B2(n5556), .A(n5557), .ZN(n5471) );
  OAI21_X2 U9183 ( .B1(n5183), .B2(n5184), .A(n5185), .ZN(n5082) );
  OAI21_X2 U9184 ( .B1(n5950), .B2(n5949), .A(n5967), .ZN(n5912) );
  OAI21_X2 U9185 ( .B1(n3734), .B2(n3735), .A(n3736), .ZN(n3558) );
  OAI21_X2 U9186 ( .B1(n4911), .B2(n4912), .A(n4913), .ZN(n4698) );
  OAI21_X2 U9187 ( .B1(n4383), .B2(n4384), .A(n4385), .ZN(n4131) );
  OAI21_X2 U9188 ( .B1(n5523), .B2(n5524), .A(n5525), .ZN(n5385) );
  OAI21_X2 U9189 ( .B1(n5155), .B2(n5156), .A(n5157), .ZN(n4970) );
  OAI21_X2 U9190 ( .B1(n3939), .B2(n3940), .A(n3941), .ZN(n3724) );
  OAI21_X2 U9191 ( .B1(n5030), .B2(n5031), .A(n5032), .ZN(n4890) );
  OAI21_X2 U9192 ( .B1(n4498), .B2(n4499), .A(n4500), .ZN(n4359) );
  OAI21_X2 U9193 ( .B1(n5596), .B2(n5597), .A(n5598), .ZN(n5511) );
  OAI21_X2 U9194 ( .B1(n5243), .B2(n5244), .A(n5245), .ZN(n5137) );
  OAI21_X2 U9195 ( .B1(n5433), .B2(n5434), .A(n5435), .ZN(n5338) );
  OAI21_X2 U9196 ( .B1(n4769), .B2(n4770), .A(n4771), .ZN(n4637) );
  OAI21_X2 U9197 ( .B1(n5036), .B2(n5037), .A(n5038), .ZN(n4896) );
  OAI21_X2 U9198 ( .B1(n4772), .B2(n4773), .A(n4774), .ZN(n4640) );
  OAI21_X2 U9199 ( .B1(n4775), .B2(n4776), .A(n4777), .ZN(n4643) );
  OAI21_X2 U9200 ( .B1(n4501), .B2(n4502), .A(n4503), .ZN(n4362) );
  OAI21_X2 U9201 ( .B1(n4504), .B2(n4505), .A(n4506), .ZN(n4365) );
  OAI21_X2 U9202 ( .B1(n4781), .B2(n4782), .A(n4783), .ZN(n4649) );
  OAI21_X2 U9203 ( .B1(n4216), .B2(n4217), .A(n4218), .ZN(n4074) );
  OAI21_X2 U9204 ( .B1(n4507), .B2(n4508), .A(n4509), .ZN(n4368) );
  OAI21_X2 U9205 ( .B1(n4219), .B2(n4220), .A(n4221), .ZN(n4077) );
  OAI21_X2 U9206 ( .B1(n4510), .B2(n4511), .A(n4512), .ZN(n4371) );
  OAI21_X2 U9207 ( .B1(n3921), .B2(n3922), .A(n3923), .ZN(n3772) );
  OAI21_X2 U9208 ( .B1(n4222), .B2(n4223), .A(n4224), .ZN(n4080) );
  OAI21_X2 U9209 ( .B1(n3924), .B2(n3925), .A(n3926), .ZN(n3775) );
  OAI21_X2 U9210 ( .B1(n4225), .B2(n4226), .A(n4227), .ZN(n4083) );
  OAI21_X2 U9211 ( .B1(n4516), .B2(n4517), .A(n4518), .ZN(n4377) );
  OAI21_X2 U9212 ( .B1(n3927), .B2(n3928), .A(n3929), .ZN(n3778) );
  OAI21_X2 U9213 ( .B1(n4228), .B2(n4229), .A(n4230), .ZN(n4086) );
  OAI21_X2 U9214 ( .B1(n3930), .B2(n3931), .A(n3932), .ZN(n3781) );
  OAI21_X2 U9215 ( .B1(n3933), .B2(n3934), .A(n3935), .ZN(n3784) );
  OAI21_X2 U9216 ( .B1(n5922), .B2(n5923), .A(n5924), .ZN(n5904) );
  OAI21_X2 U9217 ( .B1(n16381), .B2(n4065), .A(n4066), .ZN(n3911) );
  OAI21_X2 U9218 ( .B1(n5951), .B2(n2897), .A(n5937), .ZN(n5929) );
  OAI21_X2 U9219 ( .B1(n5777), .B2(n5778), .A(n5779), .ZN(n5701) );
  OAI21_X2 U9220 ( .B1(n5605), .B2(n5606), .A(n5607), .ZN(n5520) );
  OAI21_X2 U9221 ( .B1(n5704), .B2(n5705), .A(n5706), .ZN(n5560) );
  OAI21_X2 U9222 ( .B1(n5048), .B2(n5049), .A(n5050), .ZN(n4908) );
  OAI21_X2 U9223 ( .B1(n16499), .B2(n5969), .A(n5967), .ZN(n5949) );
  NOR2_X2 U9224 ( .A1(n13174), .A2(n13143), .ZN(n5969) );
  OAI21_X2 U9225 ( .B1(n16498), .B2(n5916), .A(n5896), .ZN(n5895) );
  NOR2_X2 U9226 ( .A1(n13174), .A2(n13155), .ZN(n5916) );
  OAI21_X2 U9227 ( .B1(n4790), .B2(n4791), .A(n4792), .ZN(n4658) );
  OAI21_X2 U9228 ( .B1(n4522), .B2(n4523), .A(n4524), .ZN(n4327) );
  OAI21_X2 U9229 ( .B1(n5834), .B2(n5833), .A(n5847), .ZN(n5837) );
  OAI21_X2 U9230 ( .B1(n3936), .B2(n3937), .A(n3938), .ZN(n3787) );
  OAI21_X2 U9231 ( .B1(n16473), .B2(n5135), .A(n5136), .ZN(n5027) );
  OAI21_X2 U9232 ( .B1(n16389), .B2(n4635), .A(n4636), .ZN(n4495) );
  OAI21_X2 U9233 ( .B1(n16500), .B2(n5982), .A(n5980), .ZN(n5961) );
  NOR2_X2 U9234 ( .A1(n13174), .A2(n13790), .ZN(n5982) );
  OAI21_X2 U9235 ( .B1(n3287), .B2(n3288), .A(n3197), .ZN(n3160) );
  OAI21_X2 U9236 ( .B1(n3301), .B2(n3302), .A(n3164), .ZN(n3123) );
  OAI21_X2 U9237 ( .B1(n3275), .B2(n3276), .A(n3002), .ZN(n3193) );
  OAI21_X2 U9238 ( .B1(n3281), .B2(n3282), .A(n3143), .ZN(n3148) );
  OAI21_X2 U9239 ( .B1(n3269), .B2(n3270), .A(n3176), .ZN(n3181) );
  OAI21_X2 U9240 ( .B1(n3259), .B2(n3260), .A(n2954), .ZN(n2977) );
  OAI21_X2 U9241 ( .B1(n3264), .B2(n3265), .A(n2987), .ZN(n2998) );
  OAI21_X2 U9242 ( .B1(n3412), .B2(n6003), .A(n5973), .ZN(n6002) );
  OAI21_X2 U9243 ( .B1(n2882), .B2(n6004), .A(n5979), .ZN(n5972) );
  OAI21_X2 U9244 ( .B1(n5952), .B2(n5953), .A(n5943), .ZN(n5936) );
  OAI21_X2 U9245 ( .B1(n2884), .B2(n5766), .A(n5767), .ZN(n5765) );
  OAI21_X2 U9246 ( .B1(n5736), .B2(n5737), .A(n5738), .ZN(n5735) );
  NOR2_X2 U9247 ( .A1(n5931), .A2(n5932), .ZN(n5883) );
  AOI21_X2 U9248 ( .B1(n13191), .B2(execstage_BusA[2]), .A(n16460), .ZN(n5932)
         );
  OAI21_X2 U9249 ( .B1(n5180), .B2(n5181), .A(n5182), .ZN(n5179) );
  NOR2_X2 U9250 ( .A1(n5646), .A2(n13193), .ZN(n6009) );
  OAI21_X2 U9251 ( .B1(n3255), .B2(n3256), .A(n3257), .ZN(n3254) );
  OAI21_X2 U9252 ( .B1(n5944), .B2(n5945), .A(n5954), .ZN(n5942) );
  OAI21_X2 U9253 ( .B1(n5692), .B2(n5693), .A(n5694), .ZN(n5691) );
  OAI21_X2 U9254 ( .B1(n5349), .B2(n5350), .A(n5351), .ZN(n5192) );
  OAI21_X2 U9255 ( .B1(n4092), .B2(n4093), .A(n4094), .ZN(n3827) );
  OAI21_X2 U9256 ( .B1(n5439), .B2(n5440), .A(n5441), .ZN(n5348) );
  OAI21_X2 U9257 ( .B1(n5859), .B2(n5860), .A(n5880), .ZN(n5857) );
  OAI21_X2 U9258 ( .B1(n5824), .B2(n5823), .A(n5830), .ZN(n5821) );
  OAI21_X2 U9259 ( .B1(n5552), .B2(n5553), .A(n5554), .ZN(n5551) );
  OAI21_X2 U9260 ( .B1(n5377), .B2(n5378), .A(n5379), .ZN(n5376) );
  OAI21_X2 U9261 ( .B1(n3303), .B2(n3304), .A(n3305), .ZN(n3302) );
  OAI21_X2 U9262 ( .B1(n5991), .B2(n5992), .A(n6007), .ZN(n5997) );
  OAI21_X2 U9263 ( .B1(n3790), .B2(n3791), .A(n3792), .ZN(n3472) );
  OAI21_X2 U9264 ( .B1(n4887), .B2(n4888), .A(n4889), .ZN(n4760) );
  OAI21_X2 U9265 ( .B1(n4356), .B2(n4357), .A(n4358), .ZN(n4201) );
  OAI21_X2 U9266 ( .B1(n3610), .B2(n3611), .A(n3612), .ZN(n3319) );
  OAI21_X2 U9267 ( .B1(n3613), .B2(n3614), .A(n3615), .ZN(n3353) );
  OAI21_X2 U9268 ( .B1(n3616), .B2(n3617), .A(n3618), .ZN(n3311) );
  OAI21_X2 U9269 ( .B1(n3619), .B2(n3620), .A(n3621), .ZN(n3357) );
  OAI21_X2 U9270 ( .B1(n3622), .B2(n3623), .A(n3624), .ZN(n3300) );
  OAI21_X2 U9271 ( .B1(n4213), .B2(n4214), .A(n4215), .ZN(n4073) );
  OAI21_X2 U9272 ( .B1(n4234), .B2(n4235), .A(n4236), .ZN(n4036) );
  OAI21_X2 U9273 ( .B1(n5690), .B2(n5691), .A(n5592), .ZN(n5689) );
  OAI21_X2 U9274 ( .B1(n5503), .B2(n5504), .A(n5423), .ZN(n5502) );
  OAI21_X2 U9275 ( .B1(n5236), .B2(n16485), .A(n5133), .ZN(n5235) );
  OAI21_X2 U9276 ( .B1(n5021), .B2(n5022), .A(n4886), .ZN(n5020) );
  OAI21_X2 U9277 ( .B1(n4882), .B2(n4883), .A(n4768), .ZN(n4881) );
  OAI21_X2 U9278 ( .B1(n4960), .B2(n4961), .A(n4913), .ZN(n4959) );
  OAI21_X2 U9279 ( .B1(n4688), .B2(n4689), .A(n4558), .ZN(n4687) );
  OAI21_X2 U9280 ( .B1(n4411), .B2(n4412), .A(n4385), .ZN(n4410) );
  OAI21_X2 U9281 ( .B1(n4121), .B2(n4122), .A(n4094), .ZN(n4120) );
  OAI21_X2 U9282 ( .B1(n3814), .B2(n3815), .A(n3792), .ZN(n3813) );
  OAI21_X2 U9283 ( .B1(n3457), .B2(n3458), .A(n3257), .ZN(n3456) );
  OAI21_X2 U9284 ( .B1(n5874), .B2(n5875), .A(n5876), .ZN(n5873) );
  OAI21_X2 U9285 ( .B1(n5309), .B2(n5310), .A(n5260), .ZN(n5308) );
  OAI21_X2 U9286 ( .B1(n4322), .B2(n4323), .A(n4239), .ZN(n4321) );
  OAI21_X2 U9287 ( .B1(n3719), .B2(n3720), .A(n3627), .ZN(n3718) );
  OAI21_X2 U9288 ( .B1(n16260), .B2(n3363), .A(n3364), .ZN(n3166) );
  OAI21_X2 U9289 ( .B1(n16258), .B2(n3367), .A(n3368), .ZN(n3151) );
  OAI21_X2 U9290 ( .B1(n16187), .B2(n3370), .A(n3371), .ZN(n3203) );
  OAI21_X2 U9291 ( .B1(n16262), .B2(n3360), .A(n3361), .ZN(n3027) );
  NOR2_X2 U9292 ( .A1(n4967), .A2(n5078), .ZN(n4966) );
  AOI21_X2 U9293 ( .B1(execstage_BusA[2]), .B2(n13107), .A(n5079), .ZN(n5078)
         );
  NOR2_X2 U9294 ( .A1(n4695), .A2(n4821), .ZN(n4694) );
  AOI21_X2 U9295 ( .B1(execstage_BusA[2]), .B2(n13109), .A(n4822), .ZN(n4821)
         );
  NOR2_X2 U9296 ( .A1(n5841), .A2(n16346), .ZN(n5838) );
  OAI21_X2 U9297 ( .B1(n13789), .B2(n13209), .A(n5844), .ZN(n5843) );
  NAND3_X2 U9298 ( .A1(n13795), .A2(n4957), .A3(n13109), .ZN(n4818) );
  NOR2_X2 U9299 ( .A1(n5656), .A2(n16318), .ZN(n5655) );
  OAI21_X2 U9300 ( .B1(n13150), .B2(n3565), .A(n5733), .ZN(n5732) );
  NOR2_X2 U9301 ( .A1(n5284), .A2(n16298), .ZN(n5283) );
  OAI21_X2 U9302 ( .B1(n13151), .B2(n3293), .A(n5374), .ZN(n5373) );
  OAI21_X2 U9303 ( .B1(n16405), .B2(n4758), .A(n4759), .ZN(n4756) );
  OAI21_X2 U9304 ( .B1(n4210), .B2(n4211), .A(n4212), .ZN(n4209) );
  OAI21_X2 U9305 ( .B1(n4826), .B2(n4827), .A(n4828), .ZN(n4825) );
  OAI21_X2 U9306 ( .B1(n16282), .B2(n4575), .A(n4576), .ZN(n4573) );
  OAI21_X2 U9307 ( .B1(n3551), .B2(n3552), .A(n3553), .ZN(n3550) );
  OAI21_X2 U9308 ( .B1(n16273), .B2(n4441), .A(n4442), .ZN(n4439) );
  OAI21_X2 U9309 ( .B1(n4562), .B2(n4563), .A(n4564), .ZN(n4561) );
  OAI21_X2 U9310 ( .B1(n16205), .B2(n4429), .A(n4430), .ZN(n4427) );
  OAI21_X2 U9311 ( .B1(n3538), .B2(n3539), .A(n3540), .ZN(n3537) );
  OAI21_X2 U9312 ( .B1(n16204), .B2(n4288), .A(n4289), .ZN(n4286) );
  OAI21_X2 U9313 ( .B1(n5894), .B2(n5895), .A(n5896), .ZN(n5893) );
  NAND3_X2 U9314 ( .A1(n13794), .A2(n5175), .A3(n13107), .ZN(n5075) );
  OAI21_X2 U9315 ( .B1(n8739), .B2(n13215), .A(n5405), .ZN(n5404) );
  OAI21_X2 U9316 ( .B1(n13150), .B2(n2775), .A(n5832), .ZN(n5831) );
  OAI21_X2 U9317 ( .B1(n13150), .B2(n3569), .A(n5815), .ZN(n5814) );
  OAI21_X2 U9318 ( .B1(n13789), .B2(n3555), .A(n5384), .ZN(n5383) );
  OAI21_X2 U9319 ( .B1(n2830), .B2(n13155), .A(n5678), .ZN(n5677) );
  OAI21_X2 U9320 ( .B1(n2869), .B2(n8710), .A(n5323), .ZN(n5322) );
  OAI21_X2 U9321 ( .B1(n13190), .B2(n13138), .A(n5125), .ZN(n5124) );
  OAI21_X2 U9322 ( .B1(n2775), .B2(n8710), .A(n4871), .ZN(n4870) );
  OAI21_X2 U9323 ( .B1(n13189), .B2(n13790), .A(n5928), .ZN(n5927) );
  OAI21_X2 U9324 ( .B1(n13140), .B2(n2830), .A(n5868), .ZN(n5867) );
  OAI21_X2 U9325 ( .B1(n2869), .B2(n13145), .A(n5682), .ZN(n5681) );
  OAI21_X2 U9326 ( .B1(n13140), .B2(n13212), .A(n5749), .ZN(n5748) );
  OAI21_X2 U9327 ( .B1(n13189), .B2(n13151), .A(n5940), .ZN(n5939) );
  OAI21_X2 U9328 ( .B1(n13789), .B2(n13205), .A(n5873), .ZN(n5872) );
  OAI21_X2 U9329 ( .B1(n13140), .B2(n2804), .A(n5862), .ZN(n5861) );
  OAI21_X2 U9330 ( .B1(n13153), .B2(n13215), .A(n5487), .ZN(n5486) );
  OAI21_X2 U9331 ( .B1(n5984), .B2(n5985), .A(n5986), .ZN(n5983) );
  OAI21_X2 U9332 ( .B1(n5918), .B2(n5919), .A(n5903), .ZN(n5917) );
  OAI21_X2 U9333 ( .B1(n5900), .B2(n5901), .A(n5767), .ZN(n5899) );
  INV_X4 U9334 ( .A(n13197), .ZN(n13193) );
  OAI21_X2 U9335 ( .B1(n5828), .B2(n5829), .A(n5822), .ZN(n5827) );
  OAI21_X2 U9336 ( .B1(n4556), .B2(n4557), .A(n4558), .ZN(n4555) );
  OAI21_X2 U9337 ( .B1(n16476), .B2(n5685), .A(n5686), .ZN(n5683) );
  OAI21_X2 U9338 ( .B1(n16283), .B2(n4705), .A(n4706), .ZN(n4703) );
  OAI21_X2 U9339 ( .B1(n5094), .B2(n5095), .A(n5096), .ZN(n5093) );
  OAI21_X2 U9340 ( .B1(n16272), .B2(n4300), .A(n4301), .ZN(n4298) );
  OAI21_X2 U9341 ( .B1(n3532), .B2(n3533), .A(n3534), .ZN(n3531) );
  OAI21_X2 U9342 ( .B1(n3518), .B2(n3519), .A(n3520), .ZN(n3517) );
  INV_X4 U9343 ( .A(n8809), .ZN(n13762) );
  INV_X4 U9344 ( .A(n8809), .ZN(n13761) );
  OAI21_X2 U9345 ( .B1(n5996), .B2(n5997), .A(n5998), .ZN(n5995) );
  INV_X4 U9346 ( .A(n312), .ZN(n13124) );
  INV_X4 U9347 ( .A(n312), .ZN(n13123) );
  OAI21_X2 U9348 ( .B1(n3295), .B2(n3296), .A(n3038), .ZN(n3294) );
  INV_X4 U9349 ( .A(n8809), .ZN(n13763) );
  INV_X4 U9350 ( .A(n312), .ZN(n13125) );
  AOI21_X2 U9351 ( .B1(n5836), .B2(n5835), .A(n5852), .ZN(n5834) );
  AOI21_X2 U9352 ( .B1(n5813), .B2(n5812), .A(n5816), .ZN(n5739) );
  AOI21_X2 U9353 ( .B1(n5654), .B2(n5655), .A(n5656), .ZN(n5555) );
  NOR2_X2 U9354 ( .A1(n16546), .A2(n13194), .ZN(n4797) );
  OAI21_X2 U9355 ( .B1(n3306), .B2(n3307), .A(n3116), .ZN(n3048) );
  OAI21_X2 U9356 ( .B1(n16264), .B2(n3309), .A(n3310), .ZN(n3307) );
  OAI21_X2 U9357 ( .B1(n16336), .B2(n3347), .A(n3348), .ZN(n3118) );
  OAI21_X2 U9358 ( .B1(n16325), .B2(n3351), .A(n3352), .ZN(n3110) );
  OAI21_X2 U9359 ( .B1(n16263), .B2(n3355), .A(n3356), .ZN(n3133) );
  NAND3_X2 U9360 ( .A1(n13191), .A2(n2845), .A3(n13794), .ZN(n5886) );
  OAI21_X2 U9361 ( .B1(n3141), .B2(n3142), .A(n3143), .ZN(n3138) );
  NOR2_X2 U9362 ( .A1(n5816), .A2(n16332), .ZN(n5812) );
  OAI21_X2 U9363 ( .B1(n13150), .B2(n2748), .A(n5819), .ZN(n5818) );
  NOR2_X2 U9364 ( .A1(n2998), .A2(n2999), .ZN(n2997) );
  INV_X4 U9365 ( .A(n13200), .ZN(n13194) );
  INV_X4 U9366 ( .A(n13188), .ZN(n13189) );
  INV_X4 U9367 ( .A(execstage_BusA[6]), .ZN(n13153) );
  INV_X4 U9368 ( .A(execstage_BusA[7]), .ZN(n13155) );
  INV_X4 U9369 ( .A(n8694), .ZN(n13135) );
  INV_X4 U9370 ( .A(n8648), .ZN(n13146) );
  INV_X4 U9371 ( .A(n8652), .ZN(n13141) );
  INV_X4 U9372 ( .A(execstage_BusA[5]), .ZN(n13143) );
  OAI21_X2 U9373 ( .B1(n3314), .B2(n3315), .A(n3127), .ZN(n3313) );
  INV_X4 U9374 ( .A(n8694), .ZN(n13136) );
  INV_X4 U9375 ( .A(n13188), .ZN(n13190) );
  INV_X4 U9376 ( .A(execstage_BusA[5]), .ZN(n13142) );
  INV_X4 U9377 ( .A(n8648), .ZN(n13145) );
  INV_X4 U9378 ( .A(execstage_BusA[6]), .ZN(n13154) );
  INV_X4 U9379 ( .A(execstage_BusA[5]), .ZN(n13144) );
  OAI21_X2 U9380 ( .B1(n13107), .B2(n13224), .A(n13222), .ZN(n5277) );
  NOR3_X2 U9381 ( .A1(n5543), .A2(n16457), .A3(n5544), .ZN(n5542) );
  NOR3_X2 U9382 ( .A1(n16314), .A2(n3548), .A3(n13226), .ZN(n5544) );
  AOI21_X2 U9383 ( .B1(n8649), .B2(n13165), .A(n13223), .ZN(n5546) );
  NOR3_X2 U9384 ( .A1(n16295), .A2(n16458), .A3(n5366), .ZN(n5364) );
  NOR3_X2 U9385 ( .A1(n5279), .A2(n13167), .A3(n13226), .ZN(n5366) );
  NOR2_X2 U9386 ( .A1(n13139), .A2(n3293), .ZN(n3029) );
  BUF_X4 U9387 ( .A(n13797), .Z(n12881) );
  BUF_X4 U9388 ( .A(n13797), .Z(n12882) );
  BUF_X4 U9389 ( .A(n13797), .Z(n12898) );
  BUF_X4 U9390 ( .A(n13797), .Z(n12883) );
  BUF_X4 U9391 ( .A(n13797), .Z(n12899) );
  BUF_X4 U9392 ( .A(n13797), .Z(n12884) );
  BUF_X4 U9393 ( .A(n13797), .Z(n12900) );
  BUF_X4 U9394 ( .A(n13797), .Z(n12885) );
  BUF_X4 U9395 ( .A(n13797), .Z(n12886) );
  BUF_X4 U9396 ( .A(n13797), .Z(n12901) );
  BUF_X4 U9397 ( .A(n13796), .Z(n13013) );
  BUF_X4 U9398 ( .A(n13796), .Z(n13006) );
  BUF_X4 U9399 ( .A(n13796), .Z(n13014) );
  BUF_X4 U9400 ( .A(n13796), .Z(n13007) );
  BUF_X4 U9401 ( .A(n13796), .Z(n13005) );
  INV_X4 U9402 ( .A(n13187), .ZN(n13186) );
  NOR2_X2 U9403 ( .A1(n5810), .A2(n16417), .ZN(n6023) );
  BUF_X4 U9404 ( .A(n13797), .Z(n12902) );
  BUF_X4 U9405 ( .A(n13797), .Z(n12887) );
  BUF_X4 U9406 ( .A(n13797), .Z(n12888) );
  BUF_X4 U9407 ( .A(n13797), .Z(n12903) );
  BUF_X4 U9408 ( .A(n13797), .Z(n12904) );
  BUF_X4 U9409 ( .A(n13797), .Z(n12889) );
  BUF_X4 U9410 ( .A(n13797), .Z(n12890) );
  BUF_X4 U9411 ( .A(n13797), .Z(n12905) );
  BUF_X4 U9412 ( .A(n13797), .Z(n12906) );
  BUF_X4 U9413 ( .A(n13797), .Z(n12891) );
  BUF_X4 U9414 ( .A(n13797), .Z(n12892) );
  BUF_X4 U9415 ( .A(n13797), .Z(n12907) );
  BUF_X4 U9416 ( .A(n13797), .Z(n12912) );
  BUF_X4 U9417 ( .A(n13797), .Z(n12896) );
  BUF_X4 U9418 ( .A(n13797), .Z(n12911) );
  BUF_X4 U9419 ( .A(n13797), .Z(n12895) );
  BUF_X4 U9420 ( .A(n13797), .Z(n12910) );
  BUF_X4 U9421 ( .A(n13797), .Z(n12908) );
  BUF_X4 U9422 ( .A(n13797), .Z(n12893) );
  BUF_X4 U9423 ( .A(n13797), .Z(n12894) );
  BUF_X4 U9424 ( .A(n13797), .Z(n12909) );
  BUF_X4 U9425 ( .A(n13797), .Z(n12897) );
  BUF_X4 U9426 ( .A(n13801), .Z(n10757) );
  BUF_X4 U9427 ( .A(n13801), .Z(n10748) );
  BUF_X4 U9428 ( .A(n13801), .Z(n10764) );
  BUF_X4 U9429 ( .A(n13801), .Z(n10749) );
  BUF_X4 U9430 ( .A(n13801), .Z(n10765) );
  BUF_X4 U9431 ( .A(n13801), .Z(n10750) );
  BUF_X4 U9432 ( .A(n13801), .Z(n10766) );
  BUF_X4 U9433 ( .A(n13801), .Z(n10772) );
  BUF_X4 U9434 ( .A(n13801), .Z(n10773) );
  BUF_X4 U9435 ( .A(n13801), .Z(n10758) );
  BUF_X4 U9436 ( .A(n13801), .Z(n10759) );
  BUF_X4 U9437 ( .A(n13801), .Z(n10774) );
  BUF_X4 U9438 ( .A(n13801), .Z(n10775) );
  BUF_X4 U9439 ( .A(n13801), .Z(n10753) );
  BUF_X4 U9440 ( .A(n13801), .Z(n10769) );
  BUF_X4 U9441 ( .A(n13801), .Z(n10754) );
  BUF_X4 U9442 ( .A(n13801), .Z(n10770) );
  BUF_X4 U9443 ( .A(n13801), .Z(n10755) );
  BUF_X4 U9444 ( .A(n13801), .Z(n10756) );
  BUF_X4 U9445 ( .A(n13801), .Z(n10771) );
  BUF_X4 U9446 ( .A(n13801), .Z(n10747) );
  BUF_X4 U9447 ( .A(n13801), .Z(n10762) );
  BUF_X4 U9448 ( .A(n13801), .Z(n10763) );
  BUF_X4 U9449 ( .A(n13801), .Z(n10760) );
  BUF_X4 U9450 ( .A(n13801), .Z(n10776) );
  BUF_X4 U9451 ( .A(n13801), .Z(n10746) );
  BUF_X4 U9452 ( .A(n13801), .Z(n10761) );
  BUF_X4 U9453 ( .A(n13801), .Z(n10751) );
  BUF_X4 U9454 ( .A(n13801), .Z(n10752) );
  BUF_X4 U9455 ( .A(n13801), .Z(n10767) );
  BUF_X4 U9456 ( .A(n13801), .Z(n10768) );
  BUF_X4 U9457 ( .A(n13796), .Z(n13008) );
  BUF_X4 U9458 ( .A(n13796), .Z(n13016) );
  BUF_X4 U9459 ( .A(n13796), .Z(n13009) );
  BUF_X4 U9460 ( .A(n13796), .Z(n13017) );
  BUF_X4 U9461 ( .A(n13796), .Z(n13010) );
  BUF_X4 U9462 ( .A(n13796), .Z(n13020) );
  BUF_X4 U9463 ( .A(n13796), .Z(n13012) );
  BUF_X4 U9464 ( .A(n13796), .Z(n13018) );
  BUF_X4 U9465 ( .A(n13796), .Z(n13011) );
  BUF_X4 U9466 ( .A(n13796), .Z(n13019) );
  BUF_X4 U9467 ( .A(n13796), .Z(n13015) );
  NOR2_X2 U9468 ( .A1(n2773), .A2(n16415), .ZN(n2791) );
  NOR2_X2 U9469 ( .A1(n5781), .A2(n16369), .ZN(n5796) );
  NOR2_X2 U9470 ( .A1(n2802), .A2(n16414), .ZN(n2817) );
  NOR2_X2 U9471 ( .A1(n2828), .A2(n16355), .ZN(n2840) );
  NOR2_X2 U9472 ( .A1(n6159), .A2(n6023), .ZN(n6076) );
  AOI21_X2 U9473 ( .B1(n13145), .B2(n13157), .A(n16323), .ZN(n6159) );
  INV_X4 U9474 ( .A(n13200), .ZN(n13196) );
  INV_X4 U9475 ( .A(decode_rs1_4_), .ZN(n13096) );
  AOI21_X2 U9476 ( .B1(n16539), .B2(n13194), .A(n6009), .ZN(n6018) );
  AOI222_X1 U9477 ( .A1(n4387), .A2(n16471), .B1(n4388), .B2(n8696), .C1(n3645), .C2(n8659), .ZN(n4386) );
  BUF_X4 U9478 ( .A(n13798), .Z(n10924) );
  BUF_X4 U9479 ( .A(n13798), .Z(n10942) );
  BUF_X4 U9480 ( .A(n13798), .Z(n10930) );
  BUF_X4 U9481 ( .A(n13798), .Z(n10941) );
  BUF_X4 U9482 ( .A(n13798), .Z(n10929) );
  BUF_X4 U9483 ( .A(n13798), .Z(n10936) );
  BUF_X4 U9484 ( .A(n13798), .Z(n10935) );
  BUF_X4 U9485 ( .A(n13798), .Z(n10934) );
  BUF_X4 U9486 ( .A(n13798), .Z(n10923) );
  BUF_X4 U9487 ( .A(n13798), .Z(n10938) );
  BUF_X4 U9488 ( .A(n13798), .Z(n10926) );
  BUF_X4 U9489 ( .A(n13798), .Z(n10937) );
  BUF_X4 U9490 ( .A(n13798), .Z(n10925) );
  BUF_X4 U9491 ( .A(n13798), .Z(n10932) );
  BUF_X4 U9492 ( .A(n13798), .Z(n10931) );
  BUF_X4 U9493 ( .A(n13798), .Z(n10922) );
  BUF_X4 U9494 ( .A(n13798), .Z(n10933) );
  BUF_X4 U9495 ( .A(n13798), .Z(n10940) );
  BUF_X4 U9496 ( .A(n13798), .Z(n10939) );
  BUF_X4 U9497 ( .A(n13798), .Z(n10928) );
  BUF_X4 U9498 ( .A(n13798), .Z(n10927) );
  BUF_X4 U9499 ( .A(n13798), .Z(n10921) );
  BUF_X4 U9500 ( .A(decode_rs2_1_), .Z(n10865) );
  BUF_X4 U9501 ( .A(decode_rs2_1_), .Z(n10873) );
  BUF_X4 U9502 ( .A(decode_rs2_1_), .Z(n10869) );
  BUF_X4 U9503 ( .A(decode_rs2_1_), .Z(n10877) );
  BUF_X4 U9504 ( .A(decode_rs2_1_), .Z(n10867) );
  BUF_X4 U9505 ( .A(decode_rs2_1_), .Z(n10875) );
  BUF_X4 U9506 ( .A(decode_rs2_1_), .Z(n10868) );
  BUF_X4 U9507 ( .A(decode_rs2_1_), .Z(n10876) );
  BUF_X4 U9508 ( .A(decode_rs2_1_), .Z(n10864) );
  BUF_X4 U9509 ( .A(decode_rs2_1_), .Z(n10872) );
  BUF_X4 U9510 ( .A(decode_rs2_1_), .Z(n10870) );
  BUF_X4 U9511 ( .A(decode_rs2_1_), .Z(n10878) );
  BUF_X4 U9512 ( .A(decode_rs2_1_), .Z(n10871) );
  BUF_X4 U9513 ( .A(decode_rs2_1_), .Z(n10866) );
  BUF_X4 U9514 ( .A(decode_rs2_1_), .Z(n10874) );
  BUF_X4 U9515 ( .A(decode_rs2_1_), .Z(n10863) );
  OAI21_X2 U9516 ( .B1(n16519), .B2(n5160), .A(n5161), .ZN(n3419) );
  OAI21_X2 U9517 ( .B1(n2869), .B2(n3801), .A(n5055), .ZN(n2892) );
  INV_X4 U9518 ( .A(n2873), .ZN(n16471) );
  NOR2_X2 U9519 ( .A1(n16551), .A2(n13192), .ZN(n5358) );
  OAI21_X2 U9520 ( .B1(n16520), .B2(n5160), .A(n5161), .ZN(n3395) );
  OAI21_X2 U9521 ( .B1(n16515), .B2(n5160), .A(n5266), .ZN(n4945) );
  NOR2_X2 U9522 ( .A1(n8722), .A2(n13103), .ZN(n5368) );
  OAI21_X2 U9523 ( .B1(n16517), .B2(n5160), .A(n5266), .ZN(n4944) );
  INV_X4 U9524 ( .A(n5642), .ZN(n16456) );
  INV_X4 U9525 ( .A(n5160), .ZN(n16469) );
  OAI21_X2 U9526 ( .B1(n16520), .B2(n13104), .A(n4664), .ZN(n2808) );
  OAI21_X2 U9527 ( .B1(n16515), .B2(n13104), .A(n4795), .ZN(n2831) );
  OAI21_X2 U9528 ( .B1(n13109), .B2(n13224), .A(n13222), .ZN(n5067) );
  AND2_X2 U9529 ( .A1(n13795), .A2(n8649), .ZN(n8807) );
  AOI222_X1 U9530 ( .A1(n16469), .A2(n2751), .B1(n8696), .B2(n2750), .C1(
        n16471), .C2(n2854), .ZN(n6172) );
  INV_X4 U9531 ( .A(n13200), .ZN(n13195) );
  NOR2_X2 U9532 ( .A1(n13104), .A2(n5642), .ZN(n3807) );
  OR2_X2 U9533 ( .A1(n13103), .A2(n5642), .ZN(n8808) );
  INV_X4 U9534 ( .A(n8659), .ZN(n13103) );
  INV_X4 U9535 ( .A(n8649), .ZN(n13224) );
  INV_X4 U9536 ( .A(n8649), .ZN(n13225) );
  INV_X4 U9537 ( .A(n13187), .ZN(n13185) );
  INV_X4 U9538 ( .A(n13187), .ZN(n13184) );
  INV_X4 U9539 ( .A(n13171), .ZN(n13169) );
  INV_X4 U9540 ( .A(n13171), .ZN(n13170) );
  INV_X4 U9541 ( .A(n2715), .ZN(n13223) );
  INV_X4 U9542 ( .A(n8661), .ZN(n13491) );
  INV_X4 U9543 ( .A(n8661), .ZN(n13490) );
  INV_X4 U9544 ( .A(n8699), .ZN(n13546) );
  INV_X4 U9545 ( .A(n8699), .ZN(n13545) );
  INV_X4 U9546 ( .A(n8665), .ZN(n13601) );
  INV_X4 U9547 ( .A(n8665), .ZN(n13600) );
  INV_X4 U9548 ( .A(n8666), .ZN(n13616) );
  INV_X4 U9549 ( .A(n8666), .ZN(n13615) );
  INV_X4 U9550 ( .A(n8667), .ZN(n13621) );
  INV_X4 U9551 ( .A(n8667), .ZN(n13620) );
  INV_X4 U9552 ( .A(n8700), .ZN(n13626) );
  INV_X4 U9553 ( .A(n8700), .ZN(n13625) );
  INV_X4 U9554 ( .A(n8703), .ZN(n13631) );
  INV_X4 U9555 ( .A(n8703), .ZN(n13630) );
  INV_X4 U9556 ( .A(n8704), .ZN(n13636) );
  INV_X4 U9557 ( .A(n8704), .ZN(n13635) );
  INV_X4 U9558 ( .A(n8705), .ZN(n13641) );
  INV_X4 U9559 ( .A(n8705), .ZN(n13640) );
  INV_X4 U9560 ( .A(n8706), .ZN(n13739) );
  INV_X4 U9561 ( .A(n8706), .ZN(n13738) );
  INV_X4 U9562 ( .A(n8701), .ZN(n13496) );
  INV_X4 U9563 ( .A(n8701), .ZN(n13495) );
  INV_X4 U9564 ( .A(n8702), .ZN(n13501) );
  INV_X4 U9565 ( .A(n8702), .ZN(n13500) );
  INV_X4 U9566 ( .A(n13529), .ZN(n13526) );
  INV_X4 U9567 ( .A(n13529), .ZN(n13525) );
  INV_X4 U9568 ( .A(n13534), .ZN(n13531) );
  INV_X4 U9569 ( .A(n13534), .ZN(n13530) );
  INV_X4 U9570 ( .A(n8684), .ZN(n13536) );
  INV_X4 U9571 ( .A(n8684), .ZN(n13535) );
  INV_X4 U9572 ( .A(n8685), .ZN(n13541) );
  INV_X4 U9573 ( .A(n8685), .ZN(n13540) );
  INV_X4 U9574 ( .A(n13554), .ZN(n13551) );
  INV_X4 U9575 ( .A(n13554), .ZN(n13550) );
  INV_X4 U9576 ( .A(n13559), .ZN(n13556) );
  INV_X4 U9577 ( .A(n13559), .ZN(n13555) );
  INV_X4 U9578 ( .A(n8686), .ZN(n13561) );
  INV_X4 U9579 ( .A(n8686), .ZN(n13560) );
  INV_X4 U9580 ( .A(n8687), .ZN(n13566) );
  INV_X4 U9581 ( .A(n8687), .ZN(n13565) );
  INV_X4 U9582 ( .A(n13574), .ZN(n13571) );
  INV_X4 U9583 ( .A(n13574), .ZN(n13570) );
  INV_X4 U9584 ( .A(n13579), .ZN(n13576) );
  INV_X4 U9585 ( .A(n13579), .ZN(n13575) );
  INV_X4 U9586 ( .A(n8688), .ZN(n13581) );
  INV_X4 U9587 ( .A(n8688), .ZN(n13580) );
  INV_X4 U9588 ( .A(n8689), .ZN(n13586) );
  INV_X4 U9589 ( .A(n8689), .ZN(n13585) );
  INV_X4 U9590 ( .A(n13594), .ZN(n13591) );
  INV_X4 U9591 ( .A(n13594), .ZN(n13590) );
  INV_X4 U9592 ( .A(n13599), .ZN(n13596) );
  INV_X4 U9593 ( .A(n13599), .ZN(n13595) );
  INV_X4 U9594 ( .A(n8690), .ZN(n13606) );
  INV_X4 U9595 ( .A(n8690), .ZN(n13605) );
  INV_X4 U9596 ( .A(n8691), .ZN(n13611) );
  INV_X4 U9597 ( .A(n8691), .ZN(n13610) );
  INV_X4 U9598 ( .A(n13234), .ZN(n13231) );
  INV_X4 U9599 ( .A(n13234), .ZN(n13230) );
  INV_X4 U9600 ( .A(n13289), .ZN(n13286) );
  INV_X4 U9601 ( .A(n13289), .ZN(n13285) );
  INV_X4 U9602 ( .A(n8678), .ZN(n13341) );
  INV_X4 U9603 ( .A(n8678), .ZN(n13340) );
  INV_X4 U9604 ( .A(n8681), .ZN(n13356) );
  INV_X4 U9605 ( .A(n8681), .ZN(n13355) );
  INV_X4 U9606 ( .A(n13364), .ZN(n13361) );
  INV_X4 U9607 ( .A(n13364), .ZN(n13360) );
  INV_X4 U9608 ( .A(n13369), .ZN(n13366) );
  INV_X4 U9609 ( .A(n13369), .ZN(n13365) );
  INV_X4 U9610 ( .A(n8682), .ZN(n13371) );
  INV_X4 U9611 ( .A(n8682), .ZN(n13370) );
  INV_X4 U9612 ( .A(n8683), .ZN(n13376) );
  INV_X4 U9613 ( .A(n8683), .ZN(n13375) );
  INV_X4 U9614 ( .A(n13384), .ZN(n13381) );
  INV_X4 U9615 ( .A(n13384), .ZN(n13380) );
  INV_X4 U9616 ( .A(n13482), .ZN(n13479) );
  INV_X4 U9617 ( .A(n13482), .ZN(n13478) );
  INV_X4 U9618 ( .A(n8668), .ZN(n13236) );
  INV_X4 U9619 ( .A(n8668), .ZN(n13235) );
  INV_X4 U9620 ( .A(n8669), .ZN(n13241) );
  INV_X4 U9621 ( .A(n8669), .ZN(n13240) );
  INV_X4 U9622 ( .A(n13249), .ZN(n13246) );
  INV_X4 U9623 ( .A(n13249), .ZN(n13245) );
  INV_X4 U9624 ( .A(n13254), .ZN(n13251) );
  INV_X4 U9625 ( .A(n13254), .ZN(n13250) );
  INV_X4 U9626 ( .A(n8670), .ZN(n13256) );
  INV_X4 U9627 ( .A(n8670), .ZN(n13255) );
  INV_X4 U9628 ( .A(n8671), .ZN(n13261) );
  INV_X4 U9629 ( .A(n8671), .ZN(n13260) );
  INV_X4 U9630 ( .A(n13269), .ZN(n13266) );
  INV_X4 U9631 ( .A(n13269), .ZN(n13265) );
  INV_X4 U9632 ( .A(n13274), .ZN(n13271) );
  INV_X4 U9633 ( .A(n13274), .ZN(n13270) );
  INV_X4 U9634 ( .A(n8672), .ZN(n13276) );
  INV_X4 U9635 ( .A(n8672), .ZN(n13275) );
  INV_X4 U9636 ( .A(n8673), .ZN(n13281) );
  INV_X4 U9637 ( .A(n8673), .ZN(n13280) );
  INV_X4 U9638 ( .A(n13294), .ZN(n13291) );
  INV_X4 U9639 ( .A(n13294), .ZN(n13290) );
  INV_X4 U9640 ( .A(n13299), .ZN(n13296) );
  INV_X4 U9641 ( .A(n13299), .ZN(n13295) );
  INV_X4 U9642 ( .A(n8674), .ZN(n13301) );
  INV_X4 U9643 ( .A(n8674), .ZN(n13300) );
  INV_X4 U9644 ( .A(n8675), .ZN(n13306) );
  INV_X4 U9645 ( .A(n8675), .ZN(n13305) );
  INV_X4 U9646 ( .A(n13314), .ZN(n13311) );
  INV_X4 U9647 ( .A(n13314), .ZN(n13310) );
  INV_X4 U9648 ( .A(n13319), .ZN(n13316) );
  INV_X4 U9649 ( .A(n13319), .ZN(n13315) );
  INV_X4 U9650 ( .A(n8676), .ZN(n13321) );
  INV_X4 U9651 ( .A(n8676), .ZN(n13320) );
  INV_X4 U9652 ( .A(n8677), .ZN(n13326) );
  INV_X4 U9653 ( .A(n8677), .ZN(n13325) );
  INV_X4 U9654 ( .A(n13334), .ZN(n13331) );
  INV_X4 U9655 ( .A(n13334), .ZN(n13330) );
  INV_X4 U9656 ( .A(n13339), .ZN(n13336) );
  INV_X4 U9657 ( .A(n13339), .ZN(n13335) );
  INV_X4 U9658 ( .A(n8679), .ZN(n13346) );
  INV_X4 U9659 ( .A(n8679), .ZN(n13345) );
  INV_X4 U9660 ( .A(n8680), .ZN(n13351) );
  INV_X4 U9661 ( .A(n8680), .ZN(n13350) );
  INV_X4 U9662 ( .A(n8661), .ZN(n13492) );
  INV_X4 U9663 ( .A(n8699), .ZN(n13547) );
  INV_X4 U9664 ( .A(n8665), .ZN(n13602) );
  INV_X4 U9665 ( .A(n8666), .ZN(n13617) );
  INV_X4 U9666 ( .A(n8667), .ZN(n13622) );
  INV_X4 U9667 ( .A(n8700), .ZN(n13627) );
  INV_X4 U9668 ( .A(n8703), .ZN(n13632) );
  INV_X4 U9669 ( .A(n8704), .ZN(n13637) );
  INV_X4 U9670 ( .A(n8705), .ZN(n13642) );
  INV_X4 U9671 ( .A(n8706), .ZN(n13740) );
  INV_X4 U9672 ( .A(n8701), .ZN(n13497) );
  INV_X4 U9673 ( .A(n8702), .ZN(n13502) );
  INV_X4 U9674 ( .A(n13529), .ZN(n13527) );
  INV_X4 U9675 ( .A(n13534), .ZN(n13532) );
  INV_X4 U9676 ( .A(n8684), .ZN(n13537) );
  INV_X4 U9677 ( .A(n8685), .ZN(n13542) );
  INV_X4 U9678 ( .A(n13554), .ZN(n13552) );
  INV_X4 U9679 ( .A(n13559), .ZN(n13557) );
  INV_X4 U9680 ( .A(n8686), .ZN(n13562) );
  INV_X4 U9681 ( .A(n8687), .ZN(n13567) );
  INV_X4 U9682 ( .A(n13574), .ZN(n13572) );
  INV_X4 U9683 ( .A(n13579), .ZN(n13577) );
  INV_X4 U9684 ( .A(n8688), .ZN(n13582) );
  INV_X4 U9685 ( .A(n8689), .ZN(n13587) );
  INV_X4 U9686 ( .A(n13594), .ZN(n13592) );
  INV_X4 U9687 ( .A(n13599), .ZN(n13597) );
  INV_X4 U9688 ( .A(n8690), .ZN(n13607) );
  INV_X4 U9689 ( .A(n8691), .ZN(n13612) );
  INV_X4 U9690 ( .A(n13234), .ZN(n13232) );
  INV_X4 U9691 ( .A(n13289), .ZN(n13287) );
  INV_X4 U9692 ( .A(n8678), .ZN(n13342) );
  INV_X4 U9693 ( .A(n8681), .ZN(n13357) );
  INV_X4 U9694 ( .A(n13364), .ZN(n13362) );
  INV_X4 U9695 ( .A(n13369), .ZN(n13367) );
  INV_X4 U9696 ( .A(n8682), .ZN(n13372) );
  INV_X4 U9697 ( .A(n8683), .ZN(n13377) );
  INV_X4 U9698 ( .A(n13384), .ZN(n13382) );
  INV_X4 U9699 ( .A(n13482), .ZN(n13480) );
  INV_X4 U9700 ( .A(n8668), .ZN(n13237) );
  INV_X4 U9701 ( .A(n8669), .ZN(n13242) );
  INV_X4 U9702 ( .A(n13249), .ZN(n13247) );
  INV_X4 U9703 ( .A(n13254), .ZN(n13252) );
  INV_X4 U9704 ( .A(n8670), .ZN(n13257) );
  INV_X4 U9705 ( .A(n8671), .ZN(n13262) );
  INV_X4 U9706 ( .A(n13269), .ZN(n13267) );
  INV_X4 U9707 ( .A(n13274), .ZN(n13272) );
  INV_X4 U9708 ( .A(n8672), .ZN(n13277) );
  INV_X4 U9709 ( .A(n8673), .ZN(n13282) );
  INV_X4 U9710 ( .A(n13294), .ZN(n13292) );
  INV_X4 U9711 ( .A(n13299), .ZN(n13297) );
  INV_X4 U9712 ( .A(n8674), .ZN(n13302) );
  INV_X4 U9713 ( .A(n8675), .ZN(n13307) );
  INV_X4 U9714 ( .A(n13314), .ZN(n13312) );
  INV_X4 U9715 ( .A(n13319), .ZN(n13317) );
  INV_X4 U9716 ( .A(n8676), .ZN(n13322) );
  INV_X4 U9717 ( .A(n8677), .ZN(n13327) );
  INV_X4 U9718 ( .A(n13334), .ZN(n13332) );
  INV_X4 U9719 ( .A(n13339), .ZN(n13337) );
  INV_X4 U9720 ( .A(n8679), .ZN(n13347) );
  INV_X4 U9721 ( .A(n8680), .ZN(n13352) );
  INV_X4 U9722 ( .A(n8661), .ZN(n13493) );
  INV_X4 U9723 ( .A(n8699), .ZN(n13548) );
  INV_X4 U9724 ( .A(n8665), .ZN(n13603) );
  INV_X4 U9725 ( .A(n8666), .ZN(n13618) );
  INV_X4 U9726 ( .A(n8667), .ZN(n13623) );
  INV_X4 U9727 ( .A(n8700), .ZN(n13628) );
  INV_X4 U9728 ( .A(n8703), .ZN(n13633) );
  INV_X4 U9729 ( .A(n8704), .ZN(n13638) );
  INV_X4 U9730 ( .A(n8705), .ZN(n13643) );
  INV_X4 U9731 ( .A(n8706), .ZN(n13741) );
  INV_X4 U9732 ( .A(n8701), .ZN(n13498) );
  INV_X4 U9733 ( .A(n8702), .ZN(n13503) );
  INV_X4 U9734 ( .A(n13529), .ZN(n13528) );
  INV_X4 U9735 ( .A(n13534), .ZN(n13533) );
  INV_X4 U9736 ( .A(n8684), .ZN(n13538) );
  INV_X4 U9737 ( .A(n8685), .ZN(n13543) );
  INV_X4 U9738 ( .A(n13554), .ZN(n13553) );
  INV_X4 U9739 ( .A(n13559), .ZN(n13558) );
  INV_X4 U9740 ( .A(n8686), .ZN(n13563) );
  INV_X4 U9741 ( .A(n8687), .ZN(n13568) );
  INV_X4 U9742 ( .A(n13574), .ZN(n13573) );
  INV_X4 U9743 ( .A(n13579), .ZN(n13578) );
  INV_X4 U9744 ( .A(n8688), .ZN(n13583) );
  INV_X4 U9745 ( .A(n8689), .ZN(n13588) );
  INV_X4 U9746 ( .A(n13594), .ZN(n13593) );
  INV_X4 U9747 ( .A(n13599), .ZN(n13598) );
  INV_X4 U9748 ( .A(n8690), .ZN(n13608) );
  INV_X4 U9749 ( .A(n8691), .ZN(n13613) );
  INV_X4 U9750 ( .A(n13234), .ZN(n13233) );
  INV_X4 U9751 ( .A(n13289), .ZN(n13288) );
  INV_X4 U9752 ( .A(n8678), .ZN(n13343) );
  INV_X4 U9753 ( .A(n8681), .ZN(n13358) );
  INV_X4 U9754 ( .A(n13364), .ZN(n13363) );
  INV_X4 U9755 ( .A(n13369), .ZN(n13368) );
  INV_X4 U9756 ( .A(n8682), .ZN(n13373) );
  INV_X4 U9757 ( .A(n8683), .ZN(n13378) );
  INV_X4 U9758 ( .A(n13384), .ZN(n13383) );
  INV_X4 U9759 ( .A(n13482), .ZN(n13481) );
  INV_X4 U9760 ( .A(n8668), .ZN(n13238) );
  INV_X4 U9761 ( .A(n8669), .ZN(n13243) );
  INV_X4 U9762 ( .A(n13249), .ZN(n13248) );
  INV_X4 U9763 ( .A(n13254), .ZN(n13253) );
  INV_X4 U9764 ( .A(n8670), .ZN(n13258) );
  INV_X4 U9765 ( .A(n8671), .ZN(n13263) );
  INV_X4 U9766 ( .A(n13269), .ZN(n13268) );
  INV_X4 U9767 ( .A(n13274), .ZN(n13273) );
  INV_X4 U9768 ( .A(n8672), .ZN(n13278) );
  INV_X4 U9769 ( .A(n8673), .ZN(n13283) );
  INV_X4 U9770 ( .A(n13294), .ZN(n13293) );
  INV_X4 U9771 ( .A(n13299), .ZN(n13298) );
  INV_X4 U9772 ( .A(n8674), .ZN(n13303) );
  INV_X4 U9773 ( .A(n8675), .ZN(n13308) );
  INV_X4 U9774 ( .A(n13314), .ZN(n13313) );
  INV_X4 U9775 ( .A(n13319), .ZN(n13318) );
  INV_X4 U9776 ( .A(n8676), .ZN(n13323) );
  INV_X4 U9777 ( .A(n8677), .ZN(n13328) );
  INV_X4 U9778 ( .A(n13334), .ZN(n13333) );
  INV_X4 U9779 ( .A(n13339), .ZN(n13338) );
  INV_X4 U9780 ( .A(n8679), .ZN(n13348) );
  INV_X4 U9781 ( .A(n8680), .ZN(n13353) );
  INV_X4 U9782 ( .A(n8661), .ZN(n13494) );
  INV_X4 U9783 ( .A(n8699), .ZN(n13549) );
  INV_X4 U9784 ( .A(n8665), .ZN(n13604) );
  INV_X4 U9785 ( .A(n8666), .ZN(n13619) );
  INV_X4 U9786 ( .A(n8667), .ZN(n13624) );
  INV_X4 U9787 ( .A(n8700), .ZN(n13629) );
  INV_X4 U9788 ( .A(n8703), .ZN(n13634) );
  INV_X4 U9789 ( .A(n8704), .ZN(n13639) );
  INV_X4 U9790 ( .A(n8705), .ZN(n13644) );
  INV_X4 U9791 ( .A(n8706), .ZN(n13742) );
  INV_X4 U9792 ( .A(n8701), .ZN(n13499) );
  INV_X4 U9793 ( .A(n8702), .ZN(n13504) );
  INV_X4 U9794 ( .A(n8684), .ZN(n13539) );
  INV_X4 U9795 ( .A(n8685), .ZN(n13544) );
  INV_X4 U9796 ( .A(n8686), .ZN(n13564) );
  INV_X4 U9797 ( .A(n8687), .ZN(n13569) );
  INV_X4 U9798 ( .A(n8688), .ZN(n13584) );
  INV_X4 U9799 ( .A(n8689), .ZN(n13589) );
  INV_X4 U9800 ( .A(n8690), .ZN(n13609) );
  INV_X4 U9801 ( .A(n8691), .ZN(n13614) );
  INV_X4 U9802 ( .A(n8678), .ZN(n13344) );
  INV_X4 U9803 ( .A(n8681), .ZN(n13359) );
  INV_X4 U9804 ( .A(n8682), .ZN(n13374) );
  INV_X4 U9805 ( .A(n8683), .ZN(n13379) );
  INV_X4 U9806 ( .A(n8668), .ZN(n13239) );
  INV_X4 U9807 ( .A(n8669), .ZN(n13244) );
  INV_X4 U9808 ( .A(n8670), .ZN(n13259) );
  INV_X4 U9809 ( .A(n8671), .ZN(n13264) );
  INV_X4 U9810 ( .A(n8672), .ZN(n13279) );
  INV_X4 U9811 ( .A(n8673), .ZN(n13284) );
  INV_X4 U9812 ( .A(n8674), .ZN(n13304) );
  INV_X4 U9813 ( .A(n8675), .ZN(n13309) );
  INV_X4 U9814 ( .A(n8676), .ZN(n13324) );
  INV_X4 U9815 ( .A(n8677), .ZN(n13329) );
  INV_X4 U9816 ( .A(n8679), .ZN(n13349) );
  INV_X4 U9817 ( .A(n8680), .ZN(n13354) );
  INV_X4 U9818 ( .A(n13803), .ZN(n13804) );
  INV_X4 U9819 ( .A(n13803), .ZN(n13805) );
  INV_X4 U9820 ( .A(n13803), .ZN(n13806) );
  INV_X4 U9821 ( .A(n13803), .ZN(n13807) );
  INV_X4 U9822 ( .A(n13803), .ZN(n13808) );
  AOI21_X2 U9823 ( .B1(n3883), .B2(n3884), .A(n3885), .ZN(n3734) );
  AOI21_X2 U9824 ( .B1(n3830), .B2(n3831), .A(n3832), .ZN(n3679) );
  AOI21_X2 U9825 ( .B1(n3674), .B2(n3675), .A(n3676), .ZN(n3483) );
  AOI21_X2 U9826 ( .B1(n5964), .B2(n5963), .A(n5974), .ZN(n5950) );
  AOI21_X2 U9827 ( .B1(n3819), .B2(n3820), .A(n3821), .ZN(n3669) );
  AOI21_X2 U9828 ( .B1(n4416), .B2(n4417), .A(n4418), .ZN(n4275) );
  AOI21_X2 U9829 ( .B1(n5929), .B2(n5930), .A(n5946), .ZN(n5922) );
  AOI21_X2 U9830 ( .B1(n5195), .B2(n5196), .A(n5197), .ZN(n5094) );
  AOI21_X2 U9831 ( .B1(n4327), .B2(n4328), .A(n4329), .ZN(n4234) );
  AOI21_X2 U9832 ( .B1(n3558), .B2(n3559), .A(n3560), .ZN(n3303) );
  AOI21_X2 U9833 ( .B1(n3729), .B2(n3730), .A(n3731), .ZN(n3551) );
  AOI21_X2 U9834 ( .B1(n3724), .B2(n3725), .A(n3726), .ZN(n3622) );
  AOI21_X2 U9835 ( .B1(n3714), .B2(n3715), .A(n3716), .ZN(n3538) );
  AOI21_X2 U9836 ( .B1(n4003), .B2(n4004), .A(n4005), .ZN(n3855) );
  AOI21_X2 U9837 ( .B1(n3694), .B2(n3695), .A(n3696), .ZN(n3510) );
  AOI21_X2 U9838 ( .B1(n3476), .B2(n3477), .A(n3478), .ZN(n3379) );
  AOI21_X2 U9839 ( .B1(n5027), .B2(n5028), .A(n5029), .ZN(n4887) );
  AOI21_X2 U9840 ( .B1(n3914), .B2(n3915), .A(n3916), .ZN(n3766) );
  AOI21_X2 U9841 ( .B1(n4089), .B2(n4090), .A(n4091), .ZN(n3936) );
  AOI21_X2 U9842 ( .B1(n3787), .B2(n3788), .A(n3789), .ZN(n3619) );
  AOI21_X2 U9843 ( .B1(n16504), .B2(n4931), .A(n5993), .ZN(n5991) );
  AOI21_X2 U9844 ( .B1(n4495), .B2(n4496), .A(n4497), .ZN(n4356) );
  AOI21_X2 U9845 ( .B1(n5137), .B2(n5138), .A(n5139), .ZN(n5030) );
  AOI21_X2 U9846 ( .B1(n4637), .B2(n4638), .A(n4639), .ZN(n4498) );
  AOI21_X2 U9847 ( .B1(n5695), .B2(n5696), .A(n5697), .ZN(n5596) );
  AOI21_X2 U9848 ( .B1(n5332), .B2(n5333), .A(n5334), .ZN(n5243) );
  AOI21_X2 U9849 ( .B1(n5517), .B2(n5518), .A(n5519), .ZN(n5433) );
  AOI21_X2 U9850 ( .B1(n4890), .B2(n4891), .A(n4892), .ZN(n4769) );
  AOI21_X2 U9851 ( .B1(n5143), .B2(n5144), .A(n5145), .ZN(n5036) );
  AOI21_X2 U9852 ( .B1(n4893), .B2(n4894), .A(n4895), .ZN(n4772) );
  AOI21_X2 U9853 ( .B1(n4896), .B2(n4897), .A(n4898), .ZN(n4775) );
  AOI21_X2 U9854 ( .B1(n4359), .B2(n4360), .A(n4361), .ZN(n4210) );
  AOI21_X2 U9855 ( .B1(n4640), .B2(n4641), .A(n4642), .ZN(n4501) );
  AOI21_X2 U9856 ( .B1(n4643), .B2(n4644), .A(n4645), .ZN(n4504) );
  AOI21_X2 U9857 ( .B1(n4362), .B2(n4363), .A(n4364), .ZN(n4213) );
  AOI21_X2 U9858 ( .B1(n4902), .B2(n4903), .A(n4904), .ZN(n4781) );
  AOI21_X2 U9859 ( .B1(n4646), .B2(n4647), .A(n4648), .ZN(n4507) );
  AOI21_X2 U9860 ( .B1(n4365), .B2(n4366), .A(n4367), .ZN(n4216) );
  AOI21_X2 U9861 ( .B1(n4649), .B2(n4650), .A(n4651), .ZN(n4510) );
  AOI21_X2 U9862 ( .B1(n4074), .B2(n4075), .A(n4076), .ZN(n3921) );
  AOI21_X2 U9863 ( .B1(n4368), .B2(n4369), .A(n4370), .ZN(n4219) );
  AOI21_X2 U9864 ( .B1(n3769), .B2(n3770), .A(n3771), .ZN(n3601) );
  AOI21_X2 U9865 ( .B1(n4077), .B2(n4078), .A(n4079), .ZN(n3924) );
  AOI21_X2 U9866 ( .B1(n4371), .B2(n4372), .A(n4373), .ZN(n4222) );
  AOI21_X2 U9867 ( .B1(n4655), .B2(n4656), .A(n4657), .ZN(n4516) );
  AOI21_X2 U9868 ( .B1(n4080), .B2(n4081), .A(n4082), .ZN(n3927) );
  AOI21_X2 U9869 ( .B1(n4374), .B2(n4375), .A(n4376), .ZN(n4225) );
  AOI21_X2 U9870 ( .B1(n3775), .B2(n3776), .A(n3777), .ZN(n3607) );
  AOI21_X2 U9871 ( .B1(n4083), .B2(n4084), .A(n4085), .ZN(n3930) );
  AOI21_X2 U9872 ( .B1(n4377), .B2(n4378), .A(n4379), .ZN(n4228) );
  AOI21_X2 U9873 ( .B1(n3778), .B2(n3779), .A(n3780), .ZN(n3610) );
  AOI21_X2 U9874 ( .B1(n4086), .B2(n4087), .A(n4088), .ZN(n3933) );
  AOI21_X2 U9875 ( .B1(n3781), .B2(n3782), .A(n3783), .ZN(n3613) );
  AOI21_X2 U9876 ( .B1(n3784), .B2(n3785), .A(n3786), .ZN(n3616) );
  AOI21_X2 U9877 ( .B1(n5999), .B2(n6000), .A(n5914), .ZN(n5913) );
  NOR3_X2 U9878 ( .A1(n8650), .A2(n2869), .A3(n4755), .ZN(n4639) );
  NOR3_X2 U9879 ( .A1(n3565), .A2(n13149), .A3(n5733), .ZN(n5656) );
  NOR3_X2 U9880 ( .A1(n3293), .A2(n13149), .A3(n5374), .ZN(n5284) );
  NOR3_X2 U9881 ( .A1(n8692), .A2(n13189), .A3(n5934), .ZN(n5931) );
  NOR3_X2 U9882 ( .A1(n8730), .A2(n13172), .A3(n4627), .ZN(n4497) );
  OAI21_X2 U9883 ( .B1(n13173), .B2(n8646), .A(n4488), .ZN(n4487) );
  OAI21_X2 U9884 ( .B1(n2804), .B2(n8656), .A(n3578), .ZN(n3576) );
  OAI21_X2 U9885 ( .B1(n2748), .B2(n8646), .A(n3573), .ZN(n3571) );
  OAI21_X2 U9886 ( .B1(n3569), .B2(n8730), .A(n3570), .ZN(n3568) );
  OAI21_X2 U9887 ( .B1(n13159), .B2(n8654), .A(n3567), .ZN(n3564) );
  OAI21_X2 U9888 ( .B1(n3293), .B2(n8645), .A(n3546), .ZN(n3545) );
  OAI21_X2 U9889 ( .B1(n3565), .B2(n8650), .A(n3740), .ZN(n3739) );
  OAI21_X2 U9890 ( .B1(n13173), .B2(n8647), .A(n5020), .ZN(n5019) );
  OAI21_X2 U9891 ( .B1(n13173), .B2(n8650), .A(n4881), .ZN(n4880) );
  OAI21_X2 U9892 ( .B1(n13201), .B2(n8646), .A(n4347), .ZN(n4346) );
  OAI21_X2 U9893 ( .B1(n2830), .B2(n8646), .A(n4050), .ZN(n4049) );
  OAI21_X2 U9894 ( .B1(n13149), .B2(n2830), .A(n5882), .ZN(n5881) );
  OAI21_X2 U9895 ( .B1(n2869), .B2(n8645), .A(n5127), .ZN(n5126) );
  OAI21_X2 U9896 ( .B1(n2869), .B2(n8654), .A(n4624), .ZN(n4623) );
  OAI21_X2 U9897 ( .B1(n13189), .B2(n8650), .A(n4622), .ZN(n4621) );
  OAI21_X2 U9898 ( .B1(n2830), .B2(n8647), .A(n4620), .ZN(n4619) );
  OAI21_X2 U9899 ( .B1(n13189), .B2(n8730), .A(n4345), .ZN(n4344) );
  OAI21_X2 U9900 ( .B1(n2830), .B2(n8654), .A(n4343), .ZN(n4342) );
  OAI21_X2 U9901 ( .B1(n2775), .B2(n8645), .A(n4616), .ZN(n4615) );
  OAI21_X2 U9902 ( .B1(n2804), .B2(n8650), .A(n4341), .ZN(n4340) );
  OAI21_X2 U9903 ( .B1(n2804), .B2(n13117), .A(n4048), .ZN(n4047) );
  OAI21_X2 U9904 ( .B1(n2775), .B2(n8647), .A(n4339), .ZN(n4338) );
  OAI21_X2 U9905 ( .B1(n2830), .B2(n8656), .A(n3750), .ZN(n3749) );
  OAI21_X2 U9906 ( .B1(n2775), .B2(n8654), .A(n4046), .ZN(n4045) );
  OAI21_X2 U9907 ( .B1(n2748), .B2(n8650), .A(n4044), .ZN(n4043) );
  OAI21_X2 U9908 ( .B1(n3569), .B2(n8645), .A(n4335), .ZN(n4334) );
  OAI21_X2 U9909 ( .B1(n2775), .B2(n8646), .A(n3746), .ZN(n3745) );
  OAI21_X2 U9910 ( .B1(n13157), .B2(n8647), .A(n4042), .ZN(n4041) );
  OAI21_X2 U9911 ( .B1(n2748), .B2(n13117), .A(n3744), .ZN(n3743) );
  OAI21_X2 U9912 ( .B1(n3569), .B2(n8654), .A(n3742), .ZN(n3741) );
  OAI21_X2 U9913 ( .B1(n13140), .B2(n13108), .A(n4830), .ZN(n4829) );
  OAI21_X2 U9914 ( .B1(n13150), .B2(n3145), .A(n5177), .ZN(n5176) );
  OAI21_X2 U9915 ( .B1(n13150), .B2(n13110), .A(n4959), .ZN(n4958) );
  OAI21_X2 U9916 ( .B1(n13173), .B2(n8654), .A(n4762), .ZN(n4761) );
  OAI21_X2 U9917 ( .B1(n13172), .B2(n8656), .A(n4203), .ZN(n4202) );
  OAI21_X2 U9918 ( .B1(n13793), .B2(n3293), .A(n5286), .ZN(n5285) );
  OAI21_X2 U9919 ( .B1(n13180), .B2(n8650), .A(n3563), .ZN(n3561) );
  OAI21_X2 U9920 ( .B1(n13793), .B2(n13209), .A(n5849), .ZN(n5848) );
  OAI21_X2 U9921 ( .B1(n13793), .B2(n13215), .A(n5826), .ZN(n5825) );
  OAI21_X2 U9922 ( .B1(n13793), .B2(n3565), .A(n5658), .ZN(n5657) );
  OAI21_X2 U9923 ( .B1(n13789), .B2(n13108), .A(n4969), .ZN(n4968) );
  OAI21_X2 U9924 ( .B1(n13143), .B2(n3145), .A(n4708), .ZN(n4707) );
  OAI21_X2 U9925 ( .B1(n13153), .B2(n3145), .A(n4578), .ZN(n4577) );
  OAI21_X2 U9926 ( .B1(n3555), .B2(n8647), .A(n3557), .ZN(n3554) );
  OAI21_X2 U9927 ( .B1(n8739), .B2(n3145), .A(n4444), .ZN(n4443) );
  OAI21_X2 U9928 ( .B1(n13147), .B2(n13108), .A(n4303), .ZN(n4302) );
  OAI21_X2 U9929 ( .B1(n13789), .B2(n13110), .A(n4697), .ZN(n4696) );
  OAI21_X2 U9930 ( .B1(n13140), .B2(n3201), .A(n4566), .ZN(n4565) );
  OAI21_X2 U9931 ( .B1(n13135), .B2(n3145), .A(n4012), .ZN(n4011) );
  OAI21_X2 U9932 ( .B1(n13143), .B2(n3201), .A(n4432), .ZN(n4431) );
  OAI21_X2 U9933 ( .B1(n13153), .B2(n13110), .A(n4291), .ZN(n4290) );
  OAI21_X2 U9934 ( .B1(n13137), .B2(n13108), .A(n3713), .ZN(n3712) );
  OAI21_X2 U9935 ( .B1(n8710), .B2(n13108), .A(n3536), .ZN(n3535) );
  OAI21_X2 U9936 ( .B1(n13147), .B2(n13110), .A(n4002), .ZN(n4001) );
  OAI21_X2 U9937 ( .B1(n13135), .B2(n3201), .A(n3703), .ZN(n3702) );
  OAI21_X2 U9938 ( .B1(n13141), .B2(n3201), .A(n3522), .ZN(n3521) );
  OAI21_X2 U9939 ( .B1(n13173), .B2(n8645), .A(n5235), .ZN(n5234) );
  OAI21_X2 U9940 ( .B1(n4058), .B2(n4059), .A(n3910), .ZN(n4057) );
  OAI21_X2 U9941 ( .B1(n4628), .B2(n4629), .A(n4494), .ZN(n4627) );
  OAI21_X2 U9942 ( .B1(n4267), .B2(n4268), .A(n4269), .ZN(n4126) );
  OAI21_X2 U9943 ( .B1(n3970), .B2(n3971), .A(n3972), .ZN(n3819) );
  OAI21_X2 U9944 ( .B1(n3662), .B2(n3663), .A(n3664), .ZN(n3462) );
  OAI21_X2 U9945 ( .B1(n4549), .B2(n4550), .A(n4551), .ZN(n4416) );
  OAI21_X2 U9946 ( .B1(n4193), .B2(n4194), .A(n4072), .ZN(n4071) );
  NOR2_X2 U9947 ( .A1(n13190), .A2(n8646), .ZN(n4193) );
  OAI21_X2 U9948 ( .B1(n16206), .B2(n4152), .A(n4153), .ZN(n4003) );
  OAI21_X2 U9949 ( .B1(n3855), .B2(n3856), .A(n3857), .ZN(n3704) );
  OAI21_X2 U9950 ( .B1(n16199), .B2(n4142), .A(n4143), .ZN(n3993) );
  OAI21_X2 U9951 ( .B1(n3845), .B2(n3846), .A(n3847), .ZN(n3694) );
  OAI21_X2 U9952 ( .B1(n3983), .B2(n3984), .A(n3985), .ZN(n3835) );
  OAI21_X2 U9953 ( .B1(n3684), .B2(n3685), .A(n3686), .ZN(n3496) );
  OAI21_X2 U9954 ( .B1(n3669), .B2(n3670), .A(n3671), .ZN(n3476) );
  OAI21_X2 U9955 ( .B1(n16198), .B2(n4137), .A(n4138), .ZN(n3988) );
  OAI21_X2 U9956 ( .B1(n3840), .B2(n3841), .A(n3842), .ZN(n3689) );
  OAI21_X2 U9957 ( .B1(n3978), .B2(n3979), .A(n3980), .ZN(n3830) );
  OAI21_X2 U9958 ( .B1(n3679), .B2(n3680), .A(n3681), .ZN(n3489) );
  OAI21_X2 U9959 ( .B1(n16191), .B2(n3825), .A(n3826), .ZN(n3674) );
  OAI21_X2 U9960 ( .B1(n4237), .B2(n4238), .A(n4239), .ZN(n4028) );
  OAI21_X2 U9961 ( .B1(n16373), .B2(n3918), .A(n3919), .ZN(n3769) );
  OAI21_X2 U9962 ( .B1(n5925), .B2(n2861), .A(n5876), .ZN(n5869) );
  OAI21_X2 U9963 ( .B1(n5258), .B2(n5259), .A(n5260), .ZN(n5152) );
  OAI21_X2 U9964 ( .B1(n16377), .B2(n4068), .A(n4069), .ZN(n3914) );
  OAI21_X2 U9965 ( .B1(n16497), .B2(n5898), .A(n5770), .ZN(n5769) );
  NOR2_X2 U9966 ( .A1(n13174), .A2(n13147), .ZN(n5898) );
  OAI21_X2 U9967 ( .B1(n2880), .B2(n6006), .A(n5998), .ZN(n5985) );
  OAI21_X2 U9968 ( .B1(n2885), .B2(n5920), .A(n5921), .ZN(n5919) );
  OAI21_X2 U9969 ( .B1(n3408), .B2(n6005), .A(n5986), .ZN(n5978) );
  OAI21_X2 U9970 ( .B1(n3411), .B2(n5902), .A(n5903), .ZN(n5901) );
  OAI21_X2 U9971 ( .B1(n5590), .B2(n5591), .A(n5592), .ZN(n5589) );
  NOR2_X2 U9972 ( .A1(n5142), .A2(n5225), .ZN(n5141) );
  AOI21_X2 U9973 ( .B1(n13191), .B2(n8655), .A(n5226), .ZN(n5225) );
  NOR2_X2 U9974 ( .A1(n5148), .A2(n5221), .ZN(n5147) );
  AOI21_X2 U9975 ( .B1(n13211), .B2(n8652), .A(n5222), .ZN(n5221) );
  NOR2_X2 U9976 ( .A1(n3837), .A2(n3986), .ZN(n3836) );
  AOI21_X2 U9977 ( .B1(execstage_BusA[5]), .B2(n16406), .A(n3987), .ZN(n3986)
         );
  NOR2_X2 U9978 ( .A1(n4418), .A2(n4552), .ZN(n4417) );
  AOI21_X2 U9979 ( .B1(execstage_BusA[2]), .B2(n16409), .A(n16201), .ZN(n4552)
         );
  NOR2_X2 U9980 ( .A1(n5331), .A2(n5416), .ZN(n5330) );
  AOI21_X2 U9981 ( .B1(n13176), .B2(n13120), .A(n16484), .ZN(n5416) );
  OAI21_X2 U9982 ( .B1(n4962), .B2(n4963), .A(n4964), .ZN(n4961) );
  OAI21_X2 U9983 ( .B1(n4690), .B2(n4691), .A(n4692), .ZN(n4689) );
  OAI21_X2 U9984 ( .B1(n4413), .B2(n4414), .A(n4415), .ZN(n4412) );
  OAI21_X2 U9985 ( .B1(n4123), .B2(n4124), .A(n4125), .ZN(n4122) );
  OAI21_X2 U9986 ( .B1(n3816), .B2(n3817), .A(n3818), .ZN(n3815) );
  OAI21_X2 U9987 ( .B1(n3459), .B2(n3460), .A(n3461), .ZN(n3458) );
  OAI21_X2 U9988 ( .B1(n5505), .B2(n5506), .A(n5507), .ZN(n5504) );
  OAI21_X2 U9989 ( .B1(n5421), .B2(n5422), .A(n5423), .ZN(n5420) );
  OAI21_X2 U9990 ( .B1(n4884), .B2(n4885), .A(n4886), .ZN(n4883) );
  OAI21_X2 U9991 ( .B1(n4766), .B2(n4767), .A(n4768), .ZN(n4633) );
  OAI21_X2 U9992 ( .B1(n3625), .B2(n3626), .A(n3627), .ZN(n3365) );
  OAI21_X2 U9993 ( .B1(n16181), .B2(n3262), .A(n3263), .ZN(n3260) );
  OAI21_X2 U9994 ( .B1(n16186), .B2(n3278), .A(n3279), .ZN(n3276) );
  OAI21_X2 U9995 ( .B1(n16188), .B2(n3284), .A(n3285), .ZN(n3282) );
  OAI21_X2 U9996 ( .B1(n3271), .B2(n3272), .A(n3273), .ZN(n3270) );
  OAI21_X2 U9997 ( .B1(n16184), .B2(n3267), .A(n3268), .ZN(n3265) );
  OAI21_X2 U9998 ( .B1(n16483), .B2(n5024), .A(n5025), .ZN(n5022) );
  OAI21_X2 U9999 ( .B1(n16395), .B2(n4631), .A(n4632), .ZN(n4629) );
  OAI21_X2 U10000 ( .B1(n5131), .B2(n5132), .A(n5133), .ZN(n5026) );
  OAI21_X2 U10001 ( .B1(n3763), .B2(n3764), .A(n3765), .ZN(n3589) );
  OAI21_X2 U10002 ( .B1(n3766), .B2(n3767), .A(n3768), .ZN(n3599) );
  OAI21_X2 U10003 ( .B1(n3601), .B2(n3602), .A(n3603), .ZN(n3345) );
  OAI21_X2 U10004 ( .B1(n3604), .B2(n3605), .A(n3606), .ZN(n3325) );
  OAI21_X2 U10005 ( .B1(n3607), .B2(n3608), .A(n3609), .ZN(n3349) );
  OAI21_X2 U10006 ( .B1(n3379), .B2(n3380), .A(n3381), .ZN(n2981) );
  OAI21_X2 U10007 ( .B1(n16477), .B2(n5769), .A(n5770), .ZN(n5687) );
  OAI21_X2 U10008 ( .B1(n5326), .B2(n5327), .A(n5328), .ZN(n5241) );
  OAI21_X2 U10009 ( .B1(n4350), .B2(n4351), .A(n4208), .ZN(n4349) );
  OAI21_X2 U10010 ( .B1(n3757), .B2(n3758), .A(n3594), .ZN(n3756) );
  OAI21_X2 U10011 ( .B1(n16185), .B2(n3373), .A(n3374), .ZN(n3184) );
  OAI21_X2 U10012 ( .B1(n3375), .B2(n3376), .A(n3377), .ZN(n3205) );
  OAI21_X2 U10013 ( .B1(n3386), .B2(n3387), .A(n3388), .ZN(n3219) );
  NOR2_X2 U10014 ( .A1(n5906), .A2(n5910), .ZN(n5905) );
  AOI21_X2 U10015 ( .B1(n13203), .B2(n13116), .A(n5911), .ZN(n5910) );
  NOR2_X2 U10016 ( .A1(n5513), .A2(n5583), .ZN(n5512) );
  AOI21_X2 U10017 ( .B1(n13203), .B2(n8694), .A(n5584), .ZN(n5583) );
  NOR2_X2 U10018 ( .A1(n5700), .A2(n5758), .ZN(n5699) );
  AOI21_X2 U10019 ( .B1(n13191), .B2(n13115), .A(n5759), .ZN(n5758) );
  NOR2_X2 U10020 ( .A1(n5516), .A2(n5581), .ZN(n5515) );
  AOI21_X2 U10021 ( .B1(n13191), .B2(n13118), .A(n5582), .ZN(n5581) );
  NOR2_X2 U10022 ( .A1(n5337), .A2(n5412), .ZN(n5336) );
  AOI21_X2 U10023 ( .B1(n13192), .B2(n13121), .A(n5413), .ZN(n5412) );
  NOR2_X2 U10024 ( .A1(n5340), .A2(n5410), .ZN(n5339) );
  AOI21_X2 U10025 ( .B1(n13207), .B2(n13122), .A(n5411), .ZN(n5410) );
  NOR2_X2 U10026 ( .A1(n5151), .A2(n5219), .ZN(n5150) );
  AOI21_X2 U10027 ( .B1(n13213), .B2(n8694), .A(n5220), .ZN(n5219) );
  NOR2_X2 U10028 ( .A1(n4901), .A2(n5011), .ZN(n4900) );
  AOI21_X2 U10029 ( .B1(n13211), .B2(n13120), .A(n5012), .ZN(n5011) );
  NOR2_X2 U10030 ( .A1(n5387), .A2(n5469), .ZN(n5386) );
  AOI21_X2 U10031 ( .B1(n8651), .B2(n13182), .A(n5470), .ZN(n5469) );
  NOR2_X2 U10032 ( .A1(n4907), .A2(n5007), .ZN(n4906) );
  AOI21_X2 U10033 ( .B1(n13216), .B2(n13121), .A(n5008), .ZN(n5007) );
  NOR2_X2 U10034 ( .A1(n4654), .A2(n4743), .ZN(n4653) );
  AOI21_X2 U10035 ( .B1(n13216), .B2(n8655), .A(n4744), .ZN(n4743) );
  NOR2_X2 U10036 ( .A1(n4382), .A2(n4471), .ZN(n4381) );
  AOI21_X2 U10037 ( .B1(n13160), .B2(n13120), .A(n4472), .ZN(n4471) );
  NOR2_X2 U10038 ( .A1(n4972), .A2(n5080), .ZN(n4971) );
  AOI21_X2 U10039 ( .B1(n8651), .B2(n13168), .A(n5081), .ZN(n5080) );
  NOR2_X2 U10040 ( .A1(n4700), .A2(n4823), .ZN(n4699) );
  AOI21_X2 U10041 ( .B1(n8651), .B2(n13113), .A(n4824), .ZN(n4823) );
  NOR2_X2 U10042 ( .A1(n4133), .A2(n4272), .ZN(n4132) );
  AOI21_X2 U10043 ( .B1(n8651), .B2(n16406), .A(n4273), .ZN(n4272) );
  OAI21_X2 U10044 ( .B1(n3382), .B2(n3383), .A(n3384), .ZN(n2965) );
  NOR2_X2 U10045 ( .A1(n5907), .A2(n5908), .ZN(n5870) );
  AOI21_X2 U10046 ( .B1(n13191), .B2(execstage_BusA[5]), .A(n5909), .ZN(n5908)
         );
  NOR2_X2 U10047 ( .A1(n5703), .A2(n5756), .ZN(n5702) );
  AOI21_X2 U10048 ( .B1(n13207), .B2(execstage_BusA[6]), .A(n5757), .ZN(n5756)
         );
  NOR2_X2 U10049 ( .A1(n5522), .A2(n5577), .ZN(n5521) );
  AOI21_X2 U10050 ( .B1(n13210), .B2(execstage_BusA[7]), .A(n5578), .ZN(n5577)
         );
  NOR2_X2 U10051 ( .A1(n5343), .A2(n5408), .ZN(n5342) );
  AOI21_X2 U10052 ( .B1(n13210), .B2(n13118), .A(n5409), .ZN(n5408) );
  NOR2_X2 U10053 ( .A1(n5562), .A2(n5659), .ZN(n5561) );
  AOI21_X2 U10054 ( .B1(n8651), .B2(n13158), .A(n5660), .ZN(n5659) );
  NOR2_X2 U10055 ( .A1(n5154), .A2(n5217), .ZN(n5153) );
  AOI21_X2 U10056 ( .B1(n13216), .B2(n8648), .A(n5218), .ZN(n5217) );
  NOR2_X2 U10057 ( .A1(n4910), .A2(n5005), .ZN(n4909) );
  AOI21_X2 U10058 ( .B1(n13156), .B2(n13122), .A(n5006), .ZN(n5005) );
  NOR2_X2 U10059 ( .A1(n4660), .A2(n4739), .ZN(n4659) );
  AOI21_X2 U10060 ( .B1(n13160), .B2(n8652), .A(n4740), .ZN(n4739) );
  NOR2_X2 U10061 ( .A1(n5510), .A2(n5585), .ZN(n5509) );
  AOI21_X2 U10062 ( .B1(n13176), .B2(n8652), .A(n16487), .ZN(n5585) );
  NOR2_X2 U10063 ( .A1(n4030), .A2(n4177), .ZN(n4029) );
  AOI21_X2 U10064 ( .B1(n13163), .B2(n8655), .A(n4178), .ZN(n4177) );
  NOR2_X2 U10065 ( .A1(n5306), .A2(n5398), .ZN(n5305) );
  AOI21_X2 U10066 ( .B1(execstage_BusA[6]), .B2(n13158), .A(n5399), .ZN(n5398)
         );
  NOR2_X2 U10067 ( .A1(n5202), .A2(n5297), .ZN(n5201) );
  AOI21_X2 U10068 ( .B1(execstage_BusA[5]), .B2(n13182), .A(n5298), .ZN(n5297)
         );
  NOR2_X2 U10069 ( .A1(n4020), .A2(n4169), .ZN(n4019) );
  AOI21_X2 U10070 ( .B1(n8652), .B2(n13179), .A(n4170), .ZN(n4169) );
  NOR2_X2 U10071 ( .A1(n4015), .A2(n4164), .ZN(n4014) );
  AOI21_X2 U10072 ( .B1(n13122), .B2(n13168), .A(n4165), .ZN(n4164) );
  NOR2_X2 U10073 ( .A1(n4010), .A2(n4159), .ZN(n4009) );
  AOI21_X2 U10074 ( .B1(n8648), .B2(n13107), .A(n4160), .ZN(n4159) );
  NOR2_X2 U10075 ( .A1(n3711), .A2(n3863), .ZN(n3710) );
  AOI21_X2 U10076 ( .B1(n13121), .B2(n13107), .A(n3864), .ZN(n3863) );
  NOR2_X2 U10077 ( .A1(n3706), .A2(n3858), .ZN(n3705) );
  AOI21_X2 U10078 ( .B1(n13122), .B2(n13113), .A(n3859), .ZN(n3858) );
  NOR2_X2 U10079 ( .A1(n4000), .A2(n4149), .ZN(n3999) );
  AOI21_X2 U10080 ( .B1(execstage_BusA[7]), .B2(n13109), .A(n4150), .ZN(n4149)
         );
  NOR2_X2 U10081 ( .A1(n3701), .A2(n3853), .ZN(n3700) );
  AOI21_X2 U10082 ( .B1(n8648), .B2(n13109), .A(n3854), .ZN(n3853) );
  NOR2_X2 U10083 ( .A1(n3995), .A2(n4144), .ZN(n3994) );
  AOI21_X2 U10084 ( .B1(n13116), .B2(n13112), .A(n4145), .ZN(n4144) );
  NOR2_X2 U10085 ( .A1(n3498), .A2(n3687), .ZN(n3497) );
  AOI21_X2 U10086 ( .B1(execstage_BusA[7]), .B2(n16406), .A(n3688), .ZN(n3687)
         );
  NOR2_X2 U10087 ( .A1(n5663), .A2(n5742), .ZN(n5662) );
  AOI21_X2 U10088 ( .B1(n8651), .B2(n13217), .A(n5743), .ZN(n5742) );
  NOR2_X2 U10089 ( .A1(n5473), .A2(n5558), .ZN(n5472) );
  AOI21_X2 U10090 ( .B1(n8651), .B2(n13161), .A(n5559), .ZN(n5558) );
  NOR2_X2 U10091 ( .A1(n5301), .A2(n5393), .ZN(n5300) );
  AOI21_X2 U10092 ( .B1(n13119), .B2(n13161), .A(n5394), .ZN(n5393) );
  NOR2_X2 U10093 ( .A1(n5382), .A2(n5467), .ZN(n5381) );
  AOI21_X2 U10094 ( .B1(execstage_BusA[2]), .B2(n13164), .A(n5468), .ZN(n5467)
         );
  NOR2_X2 U10095 ( .A1(n5084), .A2(n5186), .ZN(n5083) );
  AOI21_X2 U10096 ( .B1(n8651), .B2(n13179), .A(n5187), .ZN(n5186) );
  NOR2_X2 U10097 ( .A1(n3990), .A2(n4139), .ZN(n3989) );
  AOI21_X2 U10098 ( .B1(execstage_BusA[5]), .B2(n16409), .A(n4140), .ZN(n4139)
         );
  NOR2_X2 U10099 ( .A1(n3691), .A2(n3843), .ZN(n3690) );
  AOI21_X2 U10100 ( .B1(n13115), .B2(n16409), .A(n3844), .ZN(n3843) );
  NOR2_X2 U10101 ( .A1(n4128), .A2(n4270), .ZN(n4127) );
  AOI21_X2 U10102 ( .B1(execstage_BusA[2]), .B2(n13111), .A(n4271), .ZN(n4270)
         );
  NOR2_X2 U10103 ( .A1(n3491), .A2(n3682), .ZN(n3490) );
  AOI21_X2 U10104 ( .B1(execstage_BusA[6]), .B2(n13111), .A(n3683), .ZN(n3682)
         );
  NOR2_X2 U10105 ( .A1(n3464), .A2(n3665), .ZN(n3463) );
  AOI21_X2 U10106 ( .B1(execstage_BusA[2]), .B2(n16429), .A(n3666), .ZN(n3665)
         );
  NAND3_X2 U10107 ( .A1(n13794), .A2(n5072), .A3(n13113), .ZN(n4962) );
  NAND3_X2 U10108 ( .A1(n13795), .A2(n4815), .A3(n13112), .ZN(n4690) );
  NAND3_X2 U10109 ( .A1(n13795), .A2(n4546), .A3(n16406), .ZN(n4413) );
  NAND3_X2 U10110 ( .A1(n13795), .A2(n4408), .A3(n13111), .ZN(n4267) );
  NAND3_X2 U10111 ( .A1(n13795), .A2(n4264), .A3(n16431), .ZN(n4123) );
  NAND3_X2 U10112 ( .A1(n13795), .A2(n4118), .A3(n16433), .ZN(n3970) );
  NAND3_X2 U10113 ( .A1(n13795), .A2(n3967), .A3(n16435), .ZN(n3816) );
  NAND3_X2 U10114 ( .A1(n13795), .A2(n3811), .A3(n16429), .ZN(n3662) );
  NAND3_X2 U10115 ( .A1(n13795), .A2(n3659), .A3(n16427), .ZN(n3459) );
  NAND3_X2 U10116 ( .A1(n13795), .A2(n3452), .A3(n16426), .ZN(n3387) );
  OAI21_X2 U10117 ( .B1(n16382), .B2(n4199), .A(n4200), .ZN(n4197) );
  OAI21_X2 U10118 ( .B1(n16380), .B2(n3587), .A(n3588), .ZN(n3585) );
  OAI21_X2 U10119 ( .B1(n16376), .B2(n3597), .A(n3598), .ZN(n3595) );
  NAND3_X2 U10120 ( .A1(n13795), .A2(n4685), .A3(n16409), .ZN(n4549) );
  NAND3_X2 U10121 ( .A1(n13794), .A2(n3390), .A3(n16424), .ZN(n2956) );
  OAI21_X2 U10122 ( .B1(n13226), .B2(n2931), .A(n13219), .ZN(n2934) );
  OAI21_X2 U10123 ( .B1(n2869), .B2(n8647), .A(n4879), .ZN(n4878) );
  OAI21_X2 U10124 ( .B1(n13193), .B2(n13793), .A(n5646), .ZN(n6008) );
  OAI21_X2 U10125 ( .B1(n3548), .B2(n8645), .A(n3728), .ZN(n3727) );
  OAI21_X2 U10126 ( .B1(n2830), .B2(n8645), .A(n4875), .ZN(n4874) );
  NAND3_X2 U10127 ( .A1(n3223), .A2(n3224), .A3(n3225), .ZN(aluout_0[30]) );
  AOI222_X1 U10128 ( .A1(n3244), .A2(n3245), .B1(n3212), .B2(n3246), .C1(n3220), .C2(n3247), .ZN(n3224) );
  AND2_X2 U10129 ( .A1(n13808), .A2(n312), .ZN(n8809) );
  NAND3_X2 U10130 ( .A1(n16437), .A2(n13794), .A3(n3212), .ZN(n2937) );
  INV_X4 U10131 ( .A(n5264), .ZN(n13129) );
  NAND3_X2 U10132 ( .A1(n13119), .A2(n13176), .A3(n16499), .ZN(n5967) );
  NAND3_X2 U10133 ( .A1(n8651), .A2(n13176), .A3(n16500), .ZN(n5980) );
  NAND3_X2 U10134 ( .A1(execstage_BusA[7]), .A2(n13176), .A3(n16498), .ZN(
        n5896) );
  OAI21_X2 U10135 ( .B1(n4275), .B2(n4276), .A(n4277), .ZN(n4274) );
  OAI21_X2 U10136 ( .B1(n16182), .B2(n3470), .A(n3471), .ZN(n3468) );
  OAI21_X2 U10137 ( .B1(n3503), .B2(n3504), .A(n3505), .ZN(n3502) );
  OAI21_X2 U10138 ( .B1(n3483), .B2(n3484), .A(n3485), .ZN(n3482) );
  OAI21_X2 U10139 ( .B1(n4568), .B2(n4569), .A(n4570), .ZN(n4567) );
  OAI21_X2 U10140 ( .B1(n16208), .B2(n4435), .A(n4436), .ZN(n4433) );
  OAI21_X2 U10141 ( .B1(n16207), .B2(n4294), .A(n4295), .ZN(n4292) );
  OAI21_X2 U10142 ( .B1(n16202), .B2(n4423), .A(n4424), .ZN(n4421) );
  OAI21_X2 U10143 ( .B1(n16200), .B2(n4282), .A(n4283), .ZN(n4280) );
  OAI21_X2 U10144 ( .B1(n3524), .B2(n3525), .A(n3526), .ZN(n3523) );
  OAI21_X2 U10145 ( .B1(n3510), .B2(n3511), .A(n3512), .ZN(n3509) );
  INV_X4 U10146 ( .A(n2881), .ZN(n13197) );
  INV_X4 U10147 ( .A(n2881), .ZN(n13198) );
  INV_X4 U10148 ( .A(execstage_BusA[1]), .ZN(n13151) );
  INV_X4 U10149 ( .A(n2881), .ZN(n13199) );
  INV_X4 U10150 ( .A(n8692), .ZN(n13792) );
  OAI21_X2 U10151 ( .B1(n16374), .B2(n4071), .A(n4072), .ZN(n3920) );
  INV_X4 U10152 ( .A(execstage_ALUSrc), .ZN(n13787) );
  NOR2_X2 U10153 ( .A1(n8645), .A2(n13108), .ZN(n3136) );
  OAI21_X2 U10154 ( .B1(n3174), .B2(n3175), .A(n3176), .ZN(n3171) );
  NOR2_X2 U10155 ( .A1(n13174), .A2(n13793), .ZN(n3421) );
  NOR2_X2 U10156 ( .A1(n3181), .A2(n3182), .ZN(n3180) );
  OAI21_X2 U10157 ( .B1(n2985), .B2(n2986), .A(n2987), .ZN(n2982) );
  NOR3_X2 U10158 ( .A1(n8712), .A2(n2740), .A3(n2748), .ZN(n5813) );
  NOR3_X2 U10159 ( .A1(n8712), .A2(n5371), .A3(n3293), .ZN(n5282) );
  NOR3_X2 U10160 ( .A1(n8712), .A2(n2797), .A3(n2804), .ZN(n5836) );
  NOR3_X2 U10161 ( .A1(n8712), .A2(n5730), .A3(n3565), .ZN(n5654) );
  NOR3_X2 U10162 ( .A1(n2804), .A2(n13149), .A3(n5855), .ZN(n5852) );
  NOR3_X2 U10163 ( .A1(n2748), .A2(n13149), .A3(n5819), .ZN(n5816) );
  OAI21_X2 U10164 ( .B1(n13193), .B2(n8730), .A(n4764), .ZN(n4763) );
  NOR2_X2 U10165 ( .A1(n8645), .A2(n13194), .ZN(n5240) );
  OAI21_X2 U10166 ( .B1(n3327), .B2(n3328), .A(n3062), .ZN(n3083) );
  OAI21_X2 U10167 ( .B1(n3320), .B2(n3321), .A(n3065), .ZN(n3070) );
  OAI21_X2 U10168 ( .B1(n3195), .B2(n3196), .A(n3197), .ZN(n3191) );
  NOR2_X2 U10169 ( .A1(n3193), .A2(n3194), .ZN(n3192) );
  OAI21_X2 U10170 ( .B1(n16375), .B2(n3330), .A(n3331), .ZN(n3328) );
  OAI21_X2 U10171 ( .B1(n16337), .B2(n3323), .A(n3324), .ZN(n3321) );
  OAI21_X2 U10172 ( .B1(n16335), .B2(n3317), .A(n3318), .ZN(n3315) );
  OAI21_X2 U10173 ( .B1(n16379), .B2(n3340), .A(n3341), .ZN(n3089) );
  NOR2_X2 U10174 ( .A1(n13205), .A2(n13793), .ZN(n5878) );
  NAND3_X2 U10175 ( .A1(n13794), .A2(n2707), .A3(n13156), .ZN(n5736) );
  NAND3_X2 U10176 ( .A1(n13794), .A2(n5279), .A3(n13168), .ZN(n5180) );
  NOR2_X2 U10177 ( .A1(n5852), .A2(n16351), .ZN(n5835) );
  OAI21_X2 U10178 ( .B1(n13149), .B2(n13209), .A(n5855), .ZN(n5854) );
  NAND3_X2 U10179 ( .A1(n13794), .A2(n2866), .A3(n13202), .ZN(n5944) );
  NAND3_X2 U10180 ( .A1(n13794), .A2(n5547), .A3(n13163), .ZN(n5464) );
  OAI21_X2 U10181 ( .B1(n13193), .B2(n8647), .A(n16546), .ZN(n5130) );
  NAND3_X2 U10182 ( .A1(n3628), .A2(n3629), .A3(n3630), .ZN(aluout_0[28]) );
  AOI21_X2 U10183 ( .B1(n3452), .B2(n3649), .A(n16446), .ZN(n3629) );
  NOR2_X2 U10184 ( .A1(n3148), .A2(n3149), .ZN(n3147) );
  NOR2_X2 U10185 ( .A1(n16183), .A2(n2980), .ZN(n2975) );
  NOR2_X2 U10186 ( .A1(n2977), .A2(n2978), .ZN(n2976) );
  INV_X4 U10187 ( .A(n8712), .ZN(n13794) );
  INV_X4 U10188 ( .A(n13202), .ZN(n13201) );
  INV_X4 U10189 ( .A(execstage_BusA[4]), .ZN(n13140) );
  NAND3_X2 U10190 ( .A1(n13794), .A2(n16317), .A3(n13181), .ZN(n5552) );
  NAND3_X2 U10191 ( .A1(n13794), .A2(n16350), .A3(n13213), .ZN(n5824) );
  NAND3_X2 U10192 ( .A1(n13794), .A2(n16314), .A3(n13166), .ZN(n5377) );
  NAND3_X2 U10193 ( .A1(n13794), .A2(n16447), .A3(n13206), .ZN(n5859) );
  INV_X4 U10194 ( .A(n2909), .ZN(n13191) );
  INV_X4 U10195 ( .A(n13176), .ZN(n13174) );
  INV_X4 U10196 ( .A(n2909), .ZN(n13192) );
  INV_X4 U10197 ( .A(execstage_BusA[1]), .ZN(n13150) );
  INV_X4 U10198 ( .A(n13176), .ZN(n13173) );
  INV_X4 U10199 ( .A(n8651), .ZN(n13790) );
  INV_X4 U10200 ( .A(n13176), .ZN(n13172) );
  INV_X4 U10201 ( .A(execstage_BusA[8]), .ZN(n13147) );
  INV_X4 U10202 ( .A(execstage_BusA[12]), .ZN(n13137) );
  INV_X4 U10203 ( .A(execstage_BusA[16]), .ZN(n13139) );
  INV_X4 U10204 ( .A(n13206), .ZN(n13205) );
  INV_X4 U10205 ( .A(execstage_ALUSrc), .ZN(n13785) );
  INV_X4 U10206 ( .A(execstage_BusA[1]), .ZN(n13152) );
  INV_X4 U10207 ( .A(n13177), .ZN(n13175) );
  AOI222_X1 U10208 ( .A1(n3807), .A2(n3804), .B1(n16459), .B2(n2790), .C1(
        n16431), .C2(n4407), .ZN(n4400) );
  NOR2_X2 U10209 ( .A1(n8710), .A2(n3201), .ZN(n3199) );
  OAI21_X2 U10210 ( .B1(n3162), .B2(n3163), .A(n3164), .ZN(n3158) );
  NOR2_X2 U10211 ( .A1(n3160), .A2(n3161), .ZN(n3159) );
  OAI21_X2 U10212 ( .B1(n3125), .B2(n3126), .A(n3127), .ZN(n3121) );
  NOR2_X2 U10213 ( .A1(n3123), .A2(n3124), .ZN(n3122) );
  INV_X4 U10214 ( .A(n8651), .ZN(n13789) );
  INV_X4 U10215 ( .A(execstage_BusA[8]), .ZN(n13148) );
  INV_X4 U10216 ( .A(execstage_BusA[14]), .ZN(n13138) );
  INV_X4 U10217 ( .A(n13210), .ZN(n13209) );
  INV_X4 U10218 ( .A(n13213), .ZN(n13212) );
  INV_X4 U10219 ( .A(n13216), .ZN(n13215) );
  INV_X4 U10220 ( .A(execstage_ALUSrc), .ZN(n13786) );
  AOI222_X1 U10221 ( .A1(n16455), .A2(n3804), .B1(n13112), .B2(n4956), .C1(
        n3807), .C2(n4405), .ZN(n4951) );
  AOI222_X1 U10222 ( .A1(n3807), .A2(n4683), .B1(n16459), .B2(n2839), .C1(
        n16406), .C2(n4684), .ZN(n4679) );
  OAI21_X2 U10223 ( .B1(n16409), .B2(n13224), .A(n13222), .ZN(n4808) );
  NAND3_X2 U10224 ( .A1(n16474), .A2(n2869), .A3(n3808), .ZN(n4810) );
  NOR2_X2 U10225 ( .A1(n3048), .A2(n3049), .ZN(n3047) );
  NOR2_X2 U10226 ( .A1(n13804), .A2(n16156), .ZN(execstage_register_N72) );
  INV_X4 U10227 ( .A(n13181), .ZN(n13180) );
  INV_X4 U10228 ( .A(n13160), .ZN(n13159) );
  INV_X4 U10229 ( .A(n13163), .ZN(n13162) );
  INV_X4 U10230 ( .A(n13156), .ZN(n13157) );
  AOI222_X1 U10231 ( .A1(n16455), .A2(n3965), .B1(n13109), .B2(n5070), .C1(
        n3807), .C2(n5071), .ZN(n5065) );
  AOI222_X1 U10232 ( .A1(n16455), .A2(n4683), .B1(n13113), .B2(n5173), .C1(
        n3807), .C2(n5174), .ZN(n5169) );
  NOR2_X2 U10233 ( .A1(n13808), .A2(n16154), .ZN(execstage_register_N68) );
  NOR2_X2 U10234 ( .A1(n13808), .A2(n16153), .ZN(execstage_register_N69) );
  NOR2_X2 U10235 ( .A1(n13808), .A2(n16152), .ZN(execstage_register_N70) );
  NOR2_X2 U10236 ( .A1(n13808), .A2(n16157), .ZN(execstage_register_N71) );
  INV_X4 U10237 ( .A(n13168), .ZN(n13167) );
  INV_X4 U10238 ( .A(n13166), .ZN(n13165) );
  INV_X4 U10239 ( .A(n13179), .ZN(n13178) );
  OAI21_X2 U10240 ( .B1(n13163), .B2(n13224), .A(n2715), .ZN(n5647) );
  AOI222_X1 U10241 ( .A1(n16456), .A2(n2911), .B1(n2724), .B2(n4531), .C1(
        n2726), .C2(n3803), .ZN(n5362) );
  AOI222_X1 U10242 ( .A1(n16449), .A2(n2776), .B1(n13218), .B2(n5442), .C1(
        n16448), .C2(n2778), .ZN(n5363) );
  AOI222_X1 U10243 ( .A1(n16358), .A2(n16548), .B1(n5446), .B2(n13782), .C1(
        n16359), .C2(n13130), .ZN(n5361) );
  AOI222_X1 U10244 ( .A1(n16448), .A2(n2717), .B1(n5368), .B2(n3445), .C1(
        n13218), .C2(n5609), .ZN(n5541) );
  AOI222_X1 U10245 ( .A1(n16363), .A2(n16548), .B1(n5628), .B2(n13782), .C1(
        n16364), .C2(n13130), .ZN(n5539) );
  AOI222_X1 U10246 ( .A1(n16448), .A2(n2807), .B1(n5368), .B2(n3247), .C1(
        n8818), .C2(n5526), .ZN(n5454) );
  AOI222_X1 U10247 ( .A1(n16361), .A2(n16548), .B1(n5533), .B2(n13782), .C1(
        n16362), .C2(n13130), .ZN(n5452) );
  AOI222_X1 U10248 ( .A1(n16366), .A2(n16548), .B1(n5715), .B2(n13782), .C1(
        n16367), .C2(n13130), .ZN(n5634) );
  NOR3_X2 U10249 ( .A1(n5638), .A2(n16457), .A3(n5639), .ZN(n5637) );
  NOR3_X2 U10250 ( .A1(n5456), .A2(n16457), .A3(n5458), .ZN(n5455) );
  AOI21_X2 U10251 ( .B1(n8649), .B2(n13178), .A(n13223), .ZN(n5460) );
  INV_X4 U10252 ( .A(n8712), .ZN(n13795) );
  NOR2_X2 U10253 ( .A1(n13808), .A2(n16155), .ZN(execstage_register_N67) );
  NOR2_X2 U10254 ( .A1(n13808), .A2(n16170), .ZN(execstage_register_N66) );
  NOR2_X2 U10255 ( .A1(n13808), .A2(n16171), .ZN(execstage_register_N65) );
  NOR2_X2 U10256 ( .A1(n13215), .A2(n13226), .ZN(n2739) );
  OAI21_X2 U10257 ( .B1(n13217), .B2(n13225), .A(n13221), .ZN(n2742) );
  NOR2_X2 U10258 ( .A1(n13159), .A2(n13226), .ZN(n5806) );
  OAI21_X2 U10259 ( .B1(n13160), .B2(n13225), .A(n2715), .ZN(n5808) );
  NOR2_X2 U10260 ( .A1(n13180), .A2(n13226), .ZN(n5725) );
  OAI21_X2 U10261 ( .B1(n13182), .B2(n13224), .A(n2715), .ZN(n5727) );
  OAI21_X2 U10262 ( .B1(n3801), .B2(n5729), .A(n5641), .ZN(n5728) );
  AOI222_X1 U10263 ( .A1(n16323), .A2(n16548), .B1(n16456), .B2(n2732), .C1(
        n2733), .C2(n2734), .ZN(n2701) );
  AOI222_X1 U10264 ( .A1(n16449), .A2(n2717), .B1(n8648), .B2(n2713), .C1(
        n16448), .C2(n2719), .ZN(n2703) );
  AOI222_X1 U10265 ( .A1(n2723), .A2(n13783), .B1(n2724), .B2(n2725), .C1(
        n2726), .C2(n2727), .ZN(n2702) );
  AOI222_X1 U10266 ( .A1(n16548), .A2(n16330), .B1(n16458), .B2(n13202), .C1(
        n2760), .C2(n13130), .ZN(n2735) );
  AOI222_X1 U10267 ( .A1(n2724), .A2(n2749), .B1(n16448), .B2(n2750), .C1(
        n16449), .C2(n2751), .ZN(n2737) );
  AOI222_X1 U10268 ( .A1(n16456), .A2(n16465), .B1(n2726), .B2(n2753), .C1(
        n2754), .C2(n13783), .ZN(n2736) );
  AOI222_X1 U10269 ( .A1(n16456), .A2(n4104), .B1(n2726), .B2(n4668), .C1(
        n2733), .C2(n16461), .ZN(n5803) );
  AOI222_X1 U10270 ( .A1(n2724), .A2(n2805), .B1(n16448), .B2(n2806), .C1(
        n16449), .C2(n2807), .ZN(n5804) );
  AOI222_X1 U10271 ( .A1(n16417), .A2(n16548), .B1(n6022), .B2(n13782), .C1(
        n6023), .C2(n13130), .ZN(n5802) );
  AOI222_X1 U10272 ( .A1(n13114), .A2(n2706), .B1(n2707), .B2(n2708), .C1(
        n13156), .C2(n2710), .ZN(n2704) );
  OAI21_X2 U10273 ( .B1(n13158), .B2(n13224), .A(n13221), .ZN(n2708) );
  OAI21_X2 U10274 ( .B1(n13226), .B2(n2707), .A(n16321), .ZN(n2710) );
  NAND3_X2 U10275 ( .A1(n283), .A2(n163), .A3(n277), .ZN(n309) );
  INV_X4 U10276 ( .A(n8810), .ZN(n13797) );
  NOR2_X2 U10277 ( .A1(n13807), .A2(n16172), .ZN(execstage_register_N64) );
  NOR2_X2 U10278 ( .A1(n13808), .A2(n16173), .ZN(execstage_register_N63) );
  NOR2_X2 U10279 ( .A1(n13808), .A2(n16166), .ZN(execstage_register_N62) );
  NOR2_X2 U10280 ( .A1(n13807), .A2(n16167), .ZN(execstage_register_N61) );
  INV_X4 U10281 ( .A(n2919), .ZN(n13187) );
  INV_X4 U10282 ( .A(n8811), .ZN(n13796) );
  AOI21_X2 U10283 ( .B1(execstage_BusA[2]), .B2(n13173), .A(n6158), .ZN(n6150)
         );
  NOR2_X2 U10284 ( .A1(n284), .A2(n16593), .ZN(n278) );
  AOI21_X2 U10285 ( .B1(n8692), .B2(n13173), .A(n3421), .ZN(n3418) );
  NOR2_X2 U10286 ( .A1(n13205), .A2(n13226), .ZN(n2822) );
  OAI21_X2 U10287 ( .B1(n13207), .B2(n13225), .A(n13221), .ZN(n2825) );
  NOR2_X2 U10288 ( .A1(n13212), .A2(n13226), .ZN(n2766) );
  OAI21_X2 U10289 ( .B1(n13214), .B2(n13225), .A(n13221), .ZN(n2769) );
  NOR2_X2 U10290 ( .A1(n13209), .A2(n13226), .ZN(n2796) );
  OAI21_X2 U10291 ( .B1(n13211), .B2(n13225), .A(n13221), .ZN(n2799) );
  AOI222_X1 U10292 ( .A1(n16449), .A2(n2750), .B1(n13191), .B2(n2853), .C1(
        n16448), .C2(n2854), .ZN(n2843) );
  AOI222_X1 U10293 ( .A1(n2857), .A2(n13783), .B1(n2724), .B2(n2751), .C1(
        n2726), .C2(n2749), .ZN(n2842) );
  NOR3_X2 U10294 ( .A1(n3569), .A2(n13118), .A3(n6023), .ZN(n6112) );
  NOR3_X2 U10295 ( .A1(n13145), .A2(n6023), .A3(n13156), .ZN(n6149) );
  AOI211_X2 U10296 ( .C1(n16599), .C2(n16604), .A(n16605), .B(n309), .ZN(n142)
         );
  AOI211_X2 U10297 ( .C1(n2861), .C2(n2849), .A(n2760), .B(n6157), .ZN(n6116)
         );
  BUF_X4 U10298 ( .A(decode_rs1_2_), .Z(n13080) );
  BUF_X4 U10299 ( .A(decode_rs1_2_), .Z(n13068) );
  BUF_X4 U10300 ( .A(decode_rs1_2_), .Z(n13079) );
  BUF_X4 U10301 ( .A(decode_rs1_2_), .Z(n13078) );
  BUF_X4 U10302 ( .A(decode_rs1_2_), .Z(n13067) );
  BUF_X4 U10303 ( .A(decode_rs1_2_), .Z(n13066) );
  BUF_X4 U10304 ( .A(decode_rs1_2_), .Z(n13077) );
  BUF_X4 U10305 ( .A(decode_rs1_2_), .Z(n13065) );
  BUF_X4 U10306 ( .A(decode_rs1_2_), .Z(n13062) );
  BUF_X4 U10307 ( .A(decode_rs1_2_), .Z(n13074) );
  BUF_X4 U10308 ( .A(decode_rs1_2_), .Z(n13076) );
  BUF_X4 U10309 ( .A(decode_rs1_2_), .Z(n13075) );
  BUF_X4 U10310 ( .A(decode_rs1_2_), .Z(n13064) );
  BUF_X4 U10311 ( .A(decode_rs1_2_), .Z(n13063) );
  BUF_X4 U10312 ( .A(decode_rs1_2_), .Z(n13073) );
  BUF_X4 U10313 ( .A(decode_rs1_2_), .Z(n13072) );
  BUF_X4 U10314 ( .A(decode_rs1_2_), .Z(n13083) );
  BUF_X4 U10315 ( .A(decode_rs1_2_), .Z(n13071) );
  BUF_X4 U10316 ( .A(decode_rs1_2_), .Z(n13082) );
  BUF_X4 U10317 ( .A(decode_rs1_2_), .Z(n13081) );
  BUF_X4 U10318 ( .A(decode_rs1_2_), .Z(n13070) );
  BUF_X4 U10319 ( .A(decode_rs1_2_), .Z(n13069) );
  AOI222_X1 U10320 ( .A1(n16548), .A2(n16415), .B1(n13105), .B2(n2790), .C1(
        n2791), .C2(n13130), .ZN(n2762) );
  AOI222_X1 U10321 ( .A1(n2726), .A2(n2776), .B1(n16449), .B2(n2777), .C1(
        n2724), .C2(n2778), .ZN(n2764) );
  AOI222_X1 U10322 ( .A1(n16548), .A2(n16355), .B1(n13105), .B2(n2839), .C1(
        n2840), .C2(n13130), .ZN(n2818) );
  AOI222_X1 U10323 ( .A1(n2726), .A2(n2725), .B1(n16449), .B2(n2719), .C1(
        n2724), .C2(n2717), .ZN(n2820) );
  AOI222_X1 U10324 ( .A1(n16548), .A2(n16414), .B1(n13106), .B2(n2816), .C1(
        n2817), .C2(n13130), .ZN(n2792) );
  AOI222_X1 U10325 ( .A1(n2726), .A2(n2805), .B1(n16449), .B2(n2806), .C1(
        n2724), .C2(n2807), .ZN(n2794) );
  BUF_X4 U10326 ( .A(decode_rs1_2_), .Z(n13061) );
  NOR2_X2 U10327 ( .A1(n2744), .A2(n16330), .ZN(n2760) );
  NOR2_X2 U10328 ( .A1(n8652), .A2(n13182), .ZN(n5781) );
  NOR2_X2 U10329 ( .A1(n8694), .A2(n13161), .ZN(n5810) );
  NOR2_X2 U10330 ( .A1(n13119), .A2(n13207), .ZN(n2828) );
  NOR2_X2 U10331 ( .A1(n13116), .A2(n13211), .ZN(n2802) );
  NOR2_X2 U10332 ( .A1(n13115), .A2(n13214), .ZN(n2773) );
  NOR2_X2 U10333 ( .A1(n3418), .A2(n4947), .ZN(n6124) );
  AOI21_X2 U10334 ( .B1(n6152), .B2(n16329), .A(n6153), .ZN(n6151) );
  NOR2_X2 U10335 ( .A1(n3130), .A2(n13117), .ZN(n3129) );
  INV_X4 U10336 ( .A(n13719), .ZN(n13718) );
  INV_X4 U10337 ( .A(n13716), .ZN(n13715) );
  INV_X4 U10338 ( .A(n13710), .ZN(n13709) );
  INV_X4 U10339 ( .A(n13707), .ZN(n13706) );
  INV_X4 U10340 ( .A(n13704), .ZN(n13703) );
  INV_X4 U10341 ( .A(n13701), .ZN(n13700) );
  INV_X4 U10342 ( .A(n13698), .ZN(n13697) );
  INV_X4 U10343 ( .A(n13695), .ZN(n13694) );
  INV_X4 U10344 ( .A(n13692), .ZN(n13691) );
  INV_X4 U10345 ( .A(n13689), .ZN(n13688) );
  INV_X4 U10346 ( .A(n13686), .ZN(n13685) );
  INV_X4 U10347 ( .A(n13683), .ZN(n13682) );
  INV_X4 U10348 ( .A(n13677), .ZN(n13676) );
  INV_X4 U10349 ( .A(n13674), .ZN(n13673) );
  INV_X4 U10350 ( .A(n13671), .ZN(n13670) );
  INV_X4 U10351 ( .A(n13668), .ZN(n13667) );
  INV_X4 U10352 ( .A(n13665), .ZN(n13664) );
  INV_X4 U10353 ( .A(n13662), .ZN(n13661) );
  INV_X4 U10354 ( .A(n13659), .ZN(n13658) );
  INV_X4 U10355 ( .A(n13656), .ZN(n13655) );
  INV_X4 U10356 ( .A(n13653), .ZN(n13652) );
  INV_X4 U10357 ( .A(n13650), .ZN(n13649) );
  INV_X4 U10358 ( .A(n13745), .ZN(n13744) );
  INV_X4 U10359 ( .A(n13737), .ZN(n13736) );
  INV_X4 U10360 ( .A(n13734), .ZN(n13733) );
  INV_X4 U10361 ( .A(n13731), .ZN(n13730) );
  INV_X4 U10362 ( .A(n13728), .ZN(n13727) );
  INV_X4 U10363 ( .A(n13725), .ZN(n13724) );
  INV_X4 U10364 ( .A(n13722), .ZN(n13721) );
  INV_X4 U10365 ( .A(n13713), .ZN(n13712) );
  INV_X4 U10366 ( .A(n13680), .ZN(n13679) );
  INV_X4 U10367 ( .A(n13647), .ZN(n13646) );
  INV_X4 U10368 ( .A(n13719), .ZN(n13717) );
  INV_X4 U10369 ( .A(n13716), .ZN(n13714) );
  INV_X4 U10370 ( .A(n13710), .ZN(n13708) );
  INV_X4 U10371 ( .A(n13707), .ZN(n13705) );
  INV_X4 U10372 ( .A(n13704), .ZN(n13702) );
  INV_X4 U10373 ( .A(n13701), .ZN(n13699) );
  INV_X4 U10374 ( .A(n13698), .ZN(n13696) );
  INV_X4 U10375 ( .A(n13695), .ZN(n13693) );
  INV_X4 U10376 ( .A(n13692), .ZN(n13690) );
  INV_X4 U10377 ( .A(n13689), .ZN(n13687) );
  INV_X4 U10378 ( .A(n13686), .ZN(n13684) );
  INV_X4 U10379 ( .A(n13683), .ZN(n13681) );
  INV_X4 U10380 ( .A(n13677), .ZN(n13675) );
  INV_X4 U10381 ( .A(n13674), .ZN(n13672) );
  INV_X4 U10382 ( .A(n13671), .ZN(n13669) );
  INV_X4 U10383 ( .A(n13668), .ZN(n13666) );
  INV_X4 U10384 ( .A(n13665), .ZN(n13663) );
  INV_X4 U10385 ( .A(n13662), .ZN(n13660) );
  INV_X4 U10386 ( .A(n13659), .ZN(n13657) );
  INV_X4 U10387 ( .A(n13656), .ZN(n13654) );
  INV_X4 U10388 ( .A(n13653), .ZN(n13651) );
  INV_X4 U10389 ( .A(n13650), .ZN(n13648) );
  INV_X4 U10390 ( .A(n13745), .ZN(n13743) );
  INV_X4 U10391 ( .A(n13737), .ZN(n13735) );
  INV_X4 U10392 ( .A(n13734), .ZN(n13732) );
  INV_X4 U10393 ( .A(n13731), .ZN(n13729) );
  INV_X4 U10394 ( .A(n13728), .ZN(n13726) );
  INV_X4 U10395 ( .A(n13725), .ZN(n13723) );
  INV_X4 U10396 ( .A(n13722), .ZN(n13720) );
  INV_X4 U10397 ( .A(n13713), .ZN(n13711) );
  INV_X4 U10398 ( .A(n13680), .ZN(n13678) );
  INV_X4 U10399 ( .A(n13647), .ZN(n13645) );
  INV_X4 U10400 ( .A(n13459), .ZN(n13458) );
  INV_X4 U10401 ( .A(n13456), .ZN(n13455) );
  INV_X4 U10402 ( .A(n13450), .ZN(n13449) );
  INV_X4 U10403 ( .A(n13447), .ZN(n13446) );
  INV_X4 U10404 ( .A(n13444), .ZN(n13443) );
  INV_X4 U10405 ( .A(n13441), .ZN(n13440) );
  INV_X4 U10406 ( .A(n13438), .ZN(n13437) );
  INV_X4 U10407 ( .A(n13435), .ZN(n13434) );
  INV_X4 U10408 ( .A(n13432), .ZN(n13431) );
  INV_X4 U10409 ( .A(n13429), .ZN(n13428) );
  INV_X4 U10410 ( .A(n13426), .ZN(n13425) );
  INV_X4 U10411 ( .A(n13423), .ZN(n13422) );
  INV_X4 U10412 ( .A(n13417), .ZN(n13416) );
  INV_X4 U10413 ( .A(n13414), .ZN(n13413) );
  INV_X4 U10414 ( .A(n13411), .ZN(n13410) );
  INV_X4 U10415 ( .A(n13408), .ZN(n13407) );
  INV_X4 U10416 ( .A(n13405), .ZN(n13404) );
  INV_X4 U10417 ( .A(n13402), .ZN(n13401) );
  INV_X4 U10418 ( .A(n13399), .ZN(n13398) );
  INV_X4 U10419 ( .A(n13396), .ZN(n13395) );
  INV_X4 U10420 ( .A(n13393), .ZN(n13392) );
  INV_X4 U10421 ( .A(n13390), .ZN(n13389) );
  INV_X4 U10422 ( .A(n13485), .ZN(n13484) );
  INV_X4 U10423 ( .A(n13477), .ZN(n13476) );
  INV_X4 U10424 ( .A(n13474), .ZN(n13473) );
  INV_X4 U10425 ( .A(n13471), .ZN(n13470) );
  INV_X4 U10426 ( .A(n13468), .ZN(n13467) );
  INV_X4 U10427 ( .A(n13465), .ZN(n13464) );
  INV_X4 U10428 ( .A(n13462), .ZN(n13461) );
  INV_X4 U10429 ( .A(n13453), .ZN(n13452) );
  INV_X4 U10430 ( .A(n13420), .ZN(n13419) );
  INV_X4 U10431 ( .A(n13387), .ZN(n13386) );
  INV_X4 U10432 ( .A(n13459), .ZN(n13457) );
  INV_X4 U10433 ( .A(n13456), .ZN(n13454) );
  INV_X4 U10434 ( .A(n13450), .ZN(n13448) );
  INV_X4 U10435 ( .A(n13447), .ZN(n13445) );
  INV_X4 U10436 ( .A(n13444), .ZN(n13442) );
  INV_X4 U10437 ( .A(n13441), .ZN(n13439) );
  INV_X4 U10438 ( .A(n13438), .ZN(n13436) );
  INV_X4 U10439 ( .A(n13435), .ZN(n13433) );
  INV_X4 U10440 ( .A(n13432), .ZN(n13430) );
  INV_X4 U10441 ( .A(n13429), .ZN(n13427) );
  INV_X4 U10442 ( .A(n13426), .ZN(n13424) );
  INV_X4 U10443 ( .A(n13423), .ZN(n13421) );
  INV_X4 U10444 ( .A(n13417), .ZN(n13415) );
  INV_X4 U10445 ( .A(n13414), .ZN(n13412) );
  INV_X4 U10446 ( .A(n13411), .ZN(n13409) );
  INV_X4 U10447 ( .A(n13408), .ZN(n13406) );
  INV_X4 U10448 ( .A(n13405), .ZN(n13403) );
  INV_X4 U10449 ( .A(n13402), .ZN(n13400) );
  INV_X4 U10450 ( .A(n13399), .ZN(n13397) );
  INV_X4 U10451 ( .A(n13396), .ZN(n13394) );
  INV_X4 U10452 ( .A(n13393), .ZN(n13391) );
  INV_X4 U10453 ( .A(n13390), .ZN(n13388) );
  INV_X4 U10454 ( .A(n13485), .ZN(n13483) );
  INV_X4 U10455 ( .A(n13477), .ZN(n13475) );
  INV_X4 U10456 ( .A(n13474), .ZN(n13472) );
  INV_X4 U10457 ( .A(n13471), .ZN(n13469) );
  INV_X4 U10458 ( .A(n13468), .ZN(n13466) );
  INV_X4 U10459 ( .A(n13465), .ZN(n13463) );
  INV_X4 U10460 ( .A(n13462), .ZN(n13460) );
  INV_X4 U10461 ( .A(n13453), .ZN(n13451) );
  INV_X4 U10462 ( .A(n13420), .ZN(n13418) );
  INV_X4 U10463 ( .A(n13387), .ZN(n13385) );
  INV_X4 U10464 ( .A(n13802), .ZN(n13801) );
  INV_X4 U10465 ( .A(n8812), .ZN(n13747) );
  INV_X4 U10466 ( .A(n8812), .ZN(n13746) );
  INV_X4 U10467 ( .A(n8813), .ZN(n13753) );
  INV_X4 U10468 ( .A(n8813), .ZN(n13752) );
  INV_X4 U10469 ( .A(n8814), .ZN(n13750) );
  INV_X4 U10470 ( .A(n8814), .ZN(n13749) );
  INV_X4 U10471 ( .A(decode_rs1_3_), .ZN(n13095) );
  NOR2_X2 U10472 ( .A1(n13807), .A2(n16162), .ZN(execstage_register_N58) );
  NOR2_X2 U10473 ( .A1(n13807), .A2(n16160), .ZN(execstage_register_N52) );
  NOR2_X2 U10474 ( .A1(n13807), .A2(n16169), .ZN(execstage_register_N59) );
  NOR2_X2 U10475 ( .A1(n13807), .A2(n16168), .ZN(execstage_register_N60) );
  NOR2_X2 U10476 ( .A1(n13807), .A2(n16164), .ZN(execstage_register_N56) );
  NOR2_X2 U10477 ( .A1(n13807), .A2(n16165), .ZN(execstage_register_N55) );
  NOR2_X2 U10478 ( .A1(n13807), .A2(n16161), .ZN(execstage_register_N51) );
  NOR2_X2 U10479 ( .A1(n13807), .A2(n16163), .ZN(execstage_register_N57) );
  NOR2_X2 U10480 ( .A1(n13807), .A2(n16159), .ZN(execstage_register_N53) );
  NOR2_X2 U10481 ( .A1(n13807), .A2(n16158), .ZN(execstage_register_N54) );
  OAI21_X2 U10482 ( .B1(n13119), .B2(n13205), .A(n6122), .ZN(n6120) );
  NAND3_X2 U10483 ( .A1(n16354), .A2(n13140), .A3(n13191), .ZN(n6122) );
  INV_X4 U10484 ( .A(n8812), .ZN(n13748) );
  INV_X4 U10485 ( .A(n8813), .ZN(n13754) );
  INV_X4 U10486 ( .A(n8814), .ZN(n13751) );
  OAI21_X2 U10487 ( .B1(n16546), .B2(n13197), .A(n5054), .ZN(n5052) );
  NOR2_X2 U10488 ( .A1(n16521), .A2(n4797), .ZN(n5788) );
  AOI21_X2 U10489 ( .B1(n16525), .B2(n13194), .A(n4797), .ZN(n4796) );
  AOI222_X1 U10490 ( .A1(n4246), .A2(n8696), .B1(n2727), .B2(n16471), .C1(
        n2725), .C2(n8659), .ZN(n5266) );
  AOI222_X1 U10491 ( .A1(n4668), .A2(n16471), .B1(n2805), .B2(n8659), .C1(
        n4667), .C2(n8696), .ZN(n5161) );
  NAND2_X2 U10492 ( .A1(n13177), .A2(n13201), .ZN(n2873) );
  AOI222_X1 U10493 ( .A1(n3439), .A2(n8696), .B1(n3440), .B2(n16471), .C1(
        n3441), .C2(n16469), .ZN(n3438) );
  AOI222_X1 U10494 ( .A1(n16469), .A2(n2913), .B1(n16471), .B2(n2915), .C1(
        n8696), .C2(n2916), .ZN(n2912) );
  AOI222_X1 U10495 ( .A1(n13106), .A2(n16509), .B1(n13114), .B2(n2892), .C1(
        n2733), .C2(n2893), .ZN(n2863) );
  INV_X4 U10496 ( .A(n3954), .ZN(n16458) );
  NOR2_X2 U10497 ( .A1(n3434), .A2(n8712), .ZN(n4388) );
  AOI211_X2 U10498 ( .C1(n13218), .C2(n4925), .A(n4926), .B(n4927), .ZN(n4924)
         );
  AOI222_X1 U10499 ( .A1(n16516), .A2(n8649), .B1(n4947), .B2(n13130), .C1(
        n16548), .C2(n16504), .ZN(n4921) );
  AOI222_X1 U10500 ( .A1(n4935), .A2(n13783), .B1(n2724), .B2(n2719), .C1(
        n2726), .C2(n2717), .ZN(n4923) );
  AOI21_X2 U10501 ( .B1(n3398), .B2(n8807), .A(n13218), .ZN(n3399) );
  AOI21_X2 U10502 ( .B1(n8649), .B2(n13173), .A(n13223), .ZN(n3397) );
  AOI211_X2 U10503 ( .C1(n162), .C2(n163), .A(n160), .B(n13804), .ZN(
        execstage_register_N4) );
  NOR2_X2 U10504 ( .A1(n3632), .A2(n3442), .ZN(n6085) );
  AOI21_X2 U10505 ( .B1(n2866), .B2(n2867), .A(n2868), .ZN(n2865) );
  NOR3_X2 U10506 ( .A1(n4105), .A2(n3953), .A3(n16423), .ZN(n6160) );
  OAI21_X2 U10507 ( .B1(n13104), .B2(n4530), .A(n4529), .ZN(n2779) );
  OAI21_X2 U10508 ( .B1(n16427), .B2(n13225), .A(n13221), .ZN(n3797) );
  INV_X4 U10509 ( .A(n2896), .ZN(n16548) );
  OAI21_X2 U10510 ( .B1(n16435), .B2(n13225), .A(n13222), .ZN(n4110) );
  NOR3_X2 U10511 ( .A1(n16439), .A2(n13202), .A3(n3801), .ZN(n3799) );
  NOR3_X2 U10512 ( .A1(n13103), .A2(n16506), .A3(n2745), .ZN(n5639) );
  OAI21_X2 U10513 ( .B1(n16429), .B2(n13225), .A(n13222), .ZN(n3960) );
  OAI21_X2 U10514 ( .B1(n16424), .B2(n13225), .A(n13221), .ZN(n3444) );
  NOR3_X2 U10515 ( .A1(n13226), .A2(n4928), .A3(n13193), .ZN(n4927) );
  OAI21_X2 U10516 ( .B1(n16437), .B2(n13225), .A(n13221), .ZN(n3246) );
  OAI21_X2 U10517 ( .B1(n16426), .B2(n13225), .A(n13221), .ZN(n3649) );
  OAI21_X2 U10518 ( .B1(n16433), .B2(n13225), .A(n13222), .ZN(n4257) );
  OAI21_X2 U10519 ( .B1(n16431), .B2(n13224), .A(n13222), .ZN(n4402) );
  OAI21_X2 U10520 ( .B1(n13111), .B2(n13224), .A(n13222), .ZN(n4542) );
  OAI21_X2 U10521 ( .B1(n16406), .B2(n13224), .A(n13222), .ZN(n4681) );
  OAI21_X2 U10522 ( .B1(n13113), .B2(n13224), .A(n13222), .ZN(n5171) );
  OAI21_X2 U10523 ( .B1(n13112), .B2(n13224), .A(n13222), .ZN(n4953) );
  NOR2_X2 U10524 ( .A1(n13114), .A2(n2733), .ZN(n2745) );
  AOI21_X2 U10525 ( .B1(n13193), .B2(n2921), .A(n16518), .ZN(n2920) );
  AOI21_X2 U10526 ( .B1(n16404), .B2(n13194), .A(n16502), .ZN(n6013) );
  OAI21_X2 U10527 ( .B1(n13203), .B2(n13225), .A(n13221), .ZN(n2867) );
  NAND3_X2 U10528 ( .A1(n6063), .A2(n6064), .A3(n6065), .ZN(n6056) );
  NOR3_X2 U10529 ( .A1(n6073), .A2(n6074), .A3(n16322), .ZN(n6063) );
  NOR3_X2 U10530 ( .A1(n16478), .A2(n6072), .A3(n5360), .ZN(n6064) );
  NOR2_X2 U10531 ( .A1(n3806), .A2(n4114), .ZN(n4259) );
  OAI21_X2 U10532 ( .B1(n13224), .B2(n13168), .A(n13222), .ZN(n5369) );
  OAI21_X2 U10533 ( .B1(n16438), .B2(n13225), .A(n13221), .ZN(n2932) );
  NAND3_X2 U10534 ( .A1(n5643), .A2(n5644), .A3(n5645), .ZN(n4387) );
  NAND3_X2 U10535 ( .A1(n3391), .A2(n3392), .A3(n3393), .ZN(aluout_0[2]) );
  AOI222_X1 U10536 ( .A1(n3418), .A2(n13131), .B1(n2733), .B2(n3419), .C1(
        n13105), .C2(n3420), .ZN(n3392) );
  NAND3_X2 U10537 ( .A1(n142), .A2(n143), .A3(n16590), .ZN(n141) );
  NAND3_X2 U10538 ( .A1(n13113), .A2(n8647), .A3(n6103), .ZN(n6095) );
  INV_X4 U10539 ( .A(n8815), .ZN(n13764) );
  INV_X4 U10540 ( .A(n8815), .ZN(n13765) );
  INV_X4 U10541 ( .A(n2721), .ZN(n13130) );
  INV_X4 U10542 ( .A(n8816), .ZN(n13770) );
  INV_X4 U10543 ( .A(n8816), .ZN(n13771) );
  INV_X4 U10544 ( .A(n2721), .ZN(n13131) );
  INV_X4 U10545 ( .A(n8817), .ZN(n13767) );
  INV_X4 U10546 ( .A(n8817), .ZN(n13768) );
  INV_X4 U10547 ( .A(n3434), .ZN(n13171) );
  INV_X4 U10548 ( .A(n267), .ZN(n13128) );
  INV_X4 U10549 ( .A(n13799), .ZN(n13798) );
  INV_X4 U10550 ( .A(n8815), .ZN(n13766) );
  INV_X4 U10551 ( .A(n8816), .ZN(n13772) );
  INV_X4 U10552 ( .A(n8817), .ZN(n13769) );
  INV_X4 U10553 ( .A(n13219), .ZN(n13218) );
  INV_X4 U10554 ( .A(n8696), .ZN(n13104) );
  INV_X4 U10555 ( .A(n8721), .ZN(n13779) );
  INV_X4 U10556 ( .A(n8721), .ZN(n13780) );
  INV_X4 U10557 ( .A(n1236), .ZN(n13529) );
  INV_X4 U10558 ( .A(n1203), .ZN(n13534) );
  INV_X4 U10559 ( .A(n1070), .ZN(n13554) );
  INV_X4 U10560 ( .A(n1037), .ZN(n13559) );
  INV_X4 U10561 ( .A(n937), .ZN(n13574) );
  INV_X4 U10562 ( .A(n904), .ZN(n13579) );
  INV_X4 U10563 ( .A(n801), .ZN(n13594) );
  INV_X4 U10564 ( .A(n767), .ZN(n13599) );
  INV_X4 U10565 ( .A(n2575), .ZN(n13234) );
  INV_X4 U10566 ( .A(n2207), .ZN(n13289) );
  INV_X4 U10567 ( .A(n1705), .ZN(n13364) );
  INV_X4 U10568 ( .A(n1672), .ZN(n13369) );
  INV_X4 U10569 ( .A(n1572), .ZN(n13384) );
  INV_X4 U10570 ( .A(n1507), .ZN(n13482) );
  INV_X4 U10571 ( .A(n2475), .ZN(n13249) );
  INV_X4 U10572 ( .A(n2441), .ZN(n13254) );
  INV_X4 U10573 ( .A(n2340), .ZN(n13269) );
  INV_X4 U10574 ( .A(n2307), .ZN(n13274) );
  INV_X4 U10575 ( .A(n2173), .ZN(n13294) );
  INV_X4 U10576 ( .A(n2140), .ZN(n13299) );
  INV_X4 U10577 ( .A(n2040), .ZN(n13314) );
  INV_X4 U10578 ( .A(n2007), .ZN(n13319) );
  INV_X4 U10579 ( .A(n1906), .ZN(n13334) );
  INV_X4 U10580 ( .A(n1873), .ZN(n13339) );
  NAND3_X2 U10581 ( .A1(n149), .A2(n220), .A3(n160), .ZN(decode_decoder_N273)
         );
  INV_X4 U10582 ( .A(stall), .ZN(n13809) );
  AOI222_X1 U10583 ( .A1(decode_regfile_N132), .A2(n13754), .B1(n13751), .B2(
        n16559), .C1(decode_regfile_N100), .C2(n13748), .ZN(n388) );
  AOI222_X1 U10584 ( .A1(decode_regfile_N133), .A2(n13754), .B1(n13751), .B2(
        n16560), .C1(decode_regfile_N101), .C2(n13748), .ZN(n389) );
  OAI21_X2 U10585 ( .B1(n2952), .B2(n2953), .A(n2954), .ZN(n2951) );
  AOI222_X1 U10586 ( .A1(n13130), .A2(n2902), .B1(n2903), .B2(n13783), .C1(
        n16549), .C2(n16384), .ZN(n2901) );
  NOR2_X2 U10587 ( .A1(n13793), .A2(n5264), .ZN(n4931) );
  NOR2_X2 U10588 ( .A1(n13151), .A2(n5264), .ZN(n4928) );
  AOI21_X2 U10589 ( .B1(n3772), .B2(n3773), .A(n3774), .ZN(n3604) );
  AOI21_X2 U10590 ( .B1(n3911), .B2(n3912), .A(n3913), .ZN(n3763) );
  NOR2_X2 U10591 ( .A1(n13143), .A2(n2946), .ZN(n2944) );
  OAI21_X2 U10592 ( .B1(n2947), .B2(n2948), .A(n2949), .ZN(n2943) );
  AOI21_X2 U10593 ( .B1(n5975), .B2(n5976), .A(n5974), .ZN(n5963) );
  NOR3_X2 U10594 ( .A1(n3480), .A2(n8692), .A3(n3975), .ZN(n3821) );
  NOR3_X2 U10595 ( .A1(n3178), .A2(n8692), .A3(n4554), .ZN(n4418) );
  NOR3_X2 U10596 ( .A1(n8731), .A2(n13172), .A3(n4057), .ZN(n3913) );
  OAI21_X2 U10597 ( .B1(n13790), .B2(n3474), .A(n3668), .ZN(n3667) );
  OAI21_X2 U10598 ( .B1(n13173), .B2(n8653), .A(n4349), .ZN(n4348) );
  OAI21_X2 U10599 ( .B1(n13189), .B2(n8653), .A(n4052), .ZN(n4051) );
  OAI21_X2 U10600 ( .B1(n2775), .B2(n8653), .A(n3575), .ZN(n3574) );
  OAI21_X2 U10601 ( .B1(n2830), .B2(n8731), .A(n3580), .ZN(n3579) );
  OAI21_X2 U10602 ( .B1(n13172), .B2(n8733), .A(n3756), .ZN(n3755) );
  OAI21_X2 U10603 ( .B1(n2869), .B2(n8732), .A(n3754), .ZN(n3753) );
  OAI21_X2 U10604 ( .B1(n13789), .B2(n3004), .A(n3977), .ZN(n3976) );
  OAI21_X2 U10605 ( .B1(n2804), .B2(n8653), .A(n3748), .ZN(n3747) );
  OAI21_X2 U10606 ( .B1(n13172), .B2(n8732), .A(n3905), .ZN(n3904) );
  OAI21_X2 U10607 ( .B1(n13149), .B2(n3474), .A(n3969), .ZN(n3968) );
  OAI21_X2 U10608 ( .B1(n13149), .B2(n3455), .A(n3456), .ZN(n3453) );
  OAI21_X2 U10609 ( .B1(n13149), .B2(n3209), .A(n3661), .ZN(n3660) );
  OAI21_X2 U10610 ( .B1(n13149), .B2(n2946), .A(n3813), .ZN(n3812) );
  OAI21_X2 U10611 ( .B1(n2917), .B2(n3593), .A(n3594), .ZN(n3332) );
  OAI21_X2 U10612 ( .B1(n13140), .B2(n3474), .A(n3475), .ZN(n3473) );
  OAI21_X2 U10613 ( .B1(n13150), .B2(n3529), .A(n5074), .ZN(n5073) );
  OAI21_X2 U10614 ( .B1(n13150), .B2(n3515), .A(n4817), .ZN(n4816) );
  OAI21_X2 U10615 ( .B1(n13150), .B2(n3500), .A(n4548), .ZN(n4547) );
  OAI21_X2 U10616 ( .B1(n13140), .B2(n3178), .A(n4279), .ZN(n4278) );
  OAI21_X2 U10617 ( .B1(n13153), .B2(n3178), .A(n3992), .ZN(n3991) );
  OAI21_X2 U10618 ( .B1(n13147), .B2(n3178), .A(n3693), .ZN(n3692) );
  OAI21_X2 U10619 ( .B1(n13149), .B2(n3004), .A(n4266), .ZN(n4265) );
  OAI21_X2 U10620 ( .B1(n13143), .B2(n3494), .A(n3834), .ZN(n3833) );
  OAI21_X2 U10621 ( .B1(n13142), .B2(n3004), .A(n3678), .ZN(n3677) );
  OAI21_X2 U10622 ( .B1(n13150), .B2(n3178), .A(n4687), .ZN(n4686) );
  OAI21_X2 U10623 ( .B1(n13149), .B2(n3494), .A(n4410), .ZN(n4409) );
  OAI21_X2 U10624 ( .B1(n13149), .B2(n3480), .A(n4120), .ZN(n4119) );
  OAI21_X2 U10625 ( .B1(n13789), .B2(n2946), .A(n3467), .ZN(n3465) );
  OAI21_X2 U10626 ( .B1(n13172), .B2(n8713), .A(n3591), .ZN(n3590) );
  OAI21_X2 U10627 ( .B1(n13140), .B2(n3529), .A(n4702), .ZN(n4701) );
  OAI21_X2 U10628 ( .B1(n13142), .B2(n3529), .A(n4572), .ZN(n4571) );
  OAI21_X2 U10629 ( .B1(n13153), .B2(n3529), .A(n4438), .ZN(n4437) );
  OAI21_X2 U10630 ( .B1(n8739), .B2(n3529), .A(n4297), .ZN(n4296) );
  OAI21_X2 U10631 ( .B1(n13145), .B2(n3529), .A(n4007), .ZN(n4006) );
  OAI21_X2 U10632 ( .B1(n13789), .B2(n3515), .A(n4560), .ZN(n4559) );
  OAI21_X2 U10633 ( .B1(n13140), .B2(n3515), .A(n4426), .ZN(n4425) );
  OAI21_X2 U10634 ( .B1(n13142), .B2(n3515), .A(n4285), .ZN(n4284) );
  OAI21_X2 U10635 ( .B1(n13141), .B2(n3529), .A(n3708), .ZN(n3707) );
  OAI21_X2 U10636 ( .B1(n13789), .B2(n3178), .A(n4420), .ZN(n4419) );
  OAI21_X2 U10637 ( .B1(n13137), .B2(n3529), .A(n3530), .ZN(n3527) );
  OAI21_X2 U10638 ( .B1(n8739), .B2(n3515), .A(n3997), .ZN(n3996) );
  OAI21_X2 U10639 ( .B1(n13145), .B2(n3515), .A(n3698), .ZN(n3697) );
  OAI21_X2 U10640 ( .B1(n13140), .B2(n3500), .A(n4135), .ZN(n4134) );
  OAI21_X2 U10641 ( .B1(n13135), .B2(n3515), .A(n3516), .ZN(n3513) );
  OAI21_X2 U10642 ( .B1(n13153), .B2(n3500), .A(n3839), .ZN(n3838) );
  OAI21_X2 U10643 ( .B1(n13789), .B2(n3494), .A(n4130), .ZN(n4129) );
  OAI21_X2 U10644 ( .B1(n13145), .B2(n3178), .A(n3508), .ZN(n3506) );
  OAI21_X2 U10645 ( .B1(n13147), .B2(n3500), .A(n3501), .ZN(n3499) );
  OAI21_X2 U10646 ( .B1(n8739), .B2(n3494), .A(n3495), .ZN(n3492) );
  OAI21_X2 U10647 ( .B1(n13790), .B2(n3480), .A(n3823), .ZN(n3822) );
  OAI21_X2 U10648 ( .B1(n13153), .B2(n3004), .A(n3488), .ZN(n3486) );
  OAI21_X2 U10649 ( .B1(n13142), .B2(n3480), .A(n3481), .ZN(n3479) );
  OAI21_X2 U10650 ( .B1(n3581), .B2(n3582), .A(n3344), .ZN(n3343) );
  NOR2_X2 U10651 ( .A1(n2909), .A2(n8732), .ZN(n3581) );
  OAI21_X2 U10652 ( .B1(n4206), .B2(n4207), .A(n4208), .ZN(n4063) );
  OAI21_X2 U10653 ( .B1(n5989), .B2(n5990), .A(n5988), .ZN(n5959) );
  NOR2_X2 U10654 ( .A1(n13151), .A2(n13173), .ZN(n5989) );
  OAI21_X2 U10655 ( .B1(n3908), .B2(n3909), .A(n3910), .ZN(n3762) );
  OAI21_X2 U10656 ( .B1(n4492), .B2(n4493), .A(n4494), .ZN(n4355) );
  OAI21_X2 U10657 ( .B1(n16392), .B2(n3760), .A(n3761), .ZN(n3758) );
  OAI21_X2 U10658 ( .B1(n16394), .B2(n4353), .A(n4354), .ZN(n4351) );
  NOR2_X2 U10659 ( .A1(n5139), .A2(n5227), .ZN(n5138) );
  AOI21_X2 U10660 ( .B1(n13203), .B2(execstage_BusA[14]), .A(n16472), .ZN(
        n5227) );
  NOR2_X2 U10661 ( .A1(n4497), .A2(n4625), .ZN(n4496) );
  AOI21_X2 U10662 ( .B1(n13177), .B2(execstage_BusA[20]), .A(n16390), .ZN(
        n4625) );
  OAI21_X2 U10663 ( .B1(n5960), .B2(n5959), .A(n5988), .ZN(n5957) );
  NOR2_X2 U10664 ( .A1(n5334), .A2(n5414), .ZN(n5333) );
  AOI21_X2 U10665 ( .B1(n13203), .B2(execstage_BusA[12]), .A(n5415), .ZN(n5414) );
  NOR2_X2 U10666 ( .A1(n5519), .A2(n5579), .ZN(n5518) );
  AOI21_X2 U10667 ( .B1(n13207), .B2(execstage_BusA[8]), .A(n5580), .ZN(n5579)
         );
  NOR2_X2 U10668 ( .A1(n4892), .A2(n5017), .ZN(n4891) );
  AOI21_X2 U10669 ( .B1(n13203), .B2(execstage_BusA[16]), .A(n5018), .ZN(n5017) );
  NOR2_X2 U10670 ( .A1(n5145), .A2(n5223), .ZN(n5144) );
  AOI21_X2 U10671 ( .B1(n13207), .B2(execstage_BusA[12]), .A(n5224), .ZN(n5223) );
  NOR2_X2 U10672 ( .A1(n4895), .A2(n5015), .ZN(n4894) );
  AOI21_X2 U10673 ( .B1(n13192), .B2(execstage_BusA[15]), .A(n5016), .ZN(n5015) );
  NOR2_X2 U10674 ( .A1(n4898), .A2(n5013), .ZN(n4897) );
  AOI21_X2 U10675 ( .B1(n13207), .B2(execstage_BusA[14]), .A(n5014), .ZN(n5013) );
  NOR2_X2 U10676 ( .A1(n4642), .A2(n4751), .ZN(n4641) );
  AOI21_X2 U10677 ( .B1(n13192), .B2(execstage_BusA[17]), .A(n4752), .ZN(n4751) );
  NOR2_X2 U10678 ( .A1(n4361), .A2(n4485), .ZN(n4360) );
  AOI21_X2 U10679 ( .B1(n13203), .B2(execstage_BusA[20]), .A(n4486), .ZN(n4485) );
  NOR2_X2 U10680 ( .A1(n4645), .A2(n4749), .ZN(n4644) );
  AOI21_X2 U10681 ( .B1(n13207), .B2(execstage_BusA[16]), .A(n4750), .ZN(n4749) );
  NOR2_X2 U10682 ( .A1(n4364), .A2(n4483), .ZN(n4363) );
  AOI21_X2 U10683 ( .B1(n13192), .B2(execstage_BusA[19]), .A(n4484), .ZN(n4483) );
  NOR2_X2 U10684 ( .A1(n4904), .A2(n5009), .ZN(n4903) );
  AOI21_X2 U10685 ( .B1(n13213), .B2(execstage_BusA[12]), .A(n5010), .ZN(n5009) );
  NOR2_X2 U10686 ( .A1(n4648), .A2(n4747), .ZN(n4647) );
  AOI21_X2 U10687 ( .B1(n13211), .B2(execstage_BusA[15]), .A(n4748), .ZN(n4747) );
  NOR2_X2 U10688 ( .A1(n4367), .A2(n4481), .ZN(n4366) );
  AOI21_X2 U10689 ( .B1(n13206), .B2(execstage_BusA[18]), .A(n4482), .ZN(n4481) );
  NOR2_X2 U10690 ( .A1(n4651), .A2(n4745), .ZN(n4650) );
  AOI21_X2 U10691 ( .B1(n13213), .B2(execstage_BusA[14]), .A(n4746), .ZN(n4745) );
  NOR2_X2 U10692 ( .A1(n4370), .A2(n4479), .ZN(n4369) );
  AOI21_X2 U10693 ( .B1(n13210), .B2(execstage_BusA[17]), .A(n4480), .ZN(n4479) );
  NOR2_X2 U10694 ( .A1(n3771), .A2(n3900), .ZN(n3770) );
  AOI21_X2 U10695 ( .B1(n13192), .B2(execstage_BusA[23]), .A(n3901), .ZN(n3900) );
  NOR2_X2 U10696 ( .A1(n4079), .A2(n4189), .ZN(n4078) );
  AOI21_X2 U10697 ( .B1(n13210), .B2(execstage_BusA[19]), .A(n4190), .ZN(n4189) );
  NOR2_X2 U10698 ( .A1(n4373), .A2(n4477), .ZN(n4372) );
  AOI21_X2 U10699 ( .B1(n13214), .B2(execstage_BusA[16]), .A(n4478), .ZN(n4477) );
  NOR2_X2 U10700 ( .A1(n4657), .A2(n4741), .ZN(n4656) );
  AOI21_X2 U10701 ( .B1(n13158), .B2(execstage_BusA[12]), .A(n4742), .ZN(n4741) );
  NOR2_X2 U10702 ( .A1(n4082), .A2(n4187), .ZN(n4081) );
  AOI21_X2 U10703 ( .B1(n13214), .B2(execstage_BusA[18]), .A(n4188), .ZN(n4187) );
  NOR2_X2 U10704 ( .A1(n4376), .A2(n4475), .ZN(n4375) );
  AOI21_X2 U10705 ( .B1(n13216), .B2(execstage_BusA[15]), .A(n4476), .ZN(n4475) );
  NOR2_X2 U10706 ( .A1(n3777), .A2(n3896), .ZN(n3776) );
  AOI21_X2 U10707 ( .B1(n13210), .B2(execstage_BusA[21]), .A(n3897), .ZN(n3896) );
  NOR2_X2 U10708 ( .A1(n4085), .A2(n4185), .ZN(n4084) );
  AOI21_X2 U10709 ( .B1(n13217), .B2(execstage_BusA[17]), .A(n4186), .ZN(n4185) );
  NOR2_X2 U10710 ( .A1(n4379), .A2(n4473), .ZN(n4378) );
  AOI21_X2 U10711 ( .B1(n13158), .B2(execstage_BusA[14]), .A(n4474), .ZN(n4473) );
  NOR2_X2 U10712 ( .A1(n3780), .A2(n3894), .ZN(n3779) );
  AOI21_X2 U10713 ( .B1(n13214), .B2(execstage_BusA[20]), .A(n3895), .ZN(n3894) );
  NOR2_X2 U10714 ( .A1(n4088), .A2(n4183), .ZN(n4087) );
  AOI21_X2 U10715 ( .B1(n13158), .B2(execstage_BusA[16]), .A(n4184), .ZN(n4183) );
  NOR2_X2 U10716 ( .A1(n3783), .A2(n3892), .ZN(n3782) );
  AOI21_X2 U10717 ( .B1(n13216), .B2(execstage_BusA[19]), .A(n3893), .ZN(n3892) );
  NOR2_X2 U10718 ( .A1(n3786), .A2(n3890), .ZN(n3785) );
  AOI21_X2 U10719 ( .B1(n13158), .B2(execstage_BusA[18]), .A(n3891), .ZN(n3890) );
  NOR2_X2 U10720 ( .A1(n5946), .A2(n5947), .ZN(n5930) );
  AOI21_X2 U10721 ( .B1(n13203), .B2(execstage_BusA[4]), .A(n5948), .ZN(n5947)
         );
  NOR2_X2 U10722 ( .A1(n3916), .A2(n4053), .ZN(n3915) );
  AOI21_X2 U10723 ( .B1(n13203), .B2(execstage_BusA[23]), .A(n4054), .ZN(n4053) );
  NOR2_X2 U10724 ( .A1(n4091), .A2(n4181), .ZN(n4090) );
  AOI21_X2 U10725 ( .B1(n13160), .B2(execstage_BusA[15]), .A(n4182), .ZN(n4181) );
  NOR2_X2 U10726 ( .A1(n4329), .A2(n4469), .ZN(n4328) );
  AOI21_X2 U10727 ( .B1(n13181), .B2(execstage_BusA[12]), .A(n4470), .ZN(n4469) );
  NOR2_X2 U10728 ( .A1(n3789), .A2(n3888), .ZN(n3788) );
  AOI21_X2 U10729 ( .B1(n13160), .B2(execstage_BusA[17]), .A(n3889), .ZN(n3888) );
  NOR2_X2 U10730 ( .A1(n3726), .A2(n3876), .ZN(n3725) );
  AOI21_X2 U10731 ( .B1(n13166), .B2(execstage_BusA[14]), .A(n3877), .ZN(n3876) );
  NOR2_X2 U10732 ( .A1(n5697), .A2(n5760), .ZN(n5696) );
  AOI21_X2 U10733 ( .B1(n13203), .B2(execstage_BusA[8]), .A(n5761), .ZN(n5760)
         );
  NOR2_X2 U10734 ( .A1(n4076), .A2(n4191), .ZN(n4075) );
  AOI21_X2 U10735 ( .B1(n13206), .B2(execstage_BusA[20]), .A(n4192), .ZN(n4191) );
  NOR2_X2 U10736 ( .A1(n5029), .A2(n5128), .ZN(n5028) );
  AOI21_X2 U10737 ( .B1(n13177), .B2(execstage_BusA[16]), .A(n5129), .ZN(n5128) );
  NOR2_X2 U10738 ( .A1(n3731), .A2(n3881), .ZN(n3730) );
  AOI21_X2 U10739 ( .B1(n13163), .B2(execstage_BusA[15]), .A(n3882), .ZN(n3881) );
  NOR2_X2 U10740 ( .A1(n3716), .A2(n3868), .ZN(n3715) );
  AOI21_X2 U10741 ( .B1(execstage_BusA[12]), .B2(n13168), .A(n3869), .ZN(n3868) );
  NOR2_X2 U10742 ( .A1(n4005), .A2(n4154), .ZN(n4004) );
  AOI21_X2 U10743 ( .B1(execstage_BusA[8]), .B2(n13113), .A(n4155), .ZN(n4154)
         );
  NOR2_X2 U10744 ( .A1(n3696), .A2(n3848), .ZN(n3695) );
  AOI21_X2 U10745 ( .B1(execstage_BusA[8]), .B2(n13112), .A(n3849), .ZN(n3848)
         );
  NOR2_X2 U10746 ( .A1(n5197), .A2(n5292), .ZN(n5196) );
  AOI21_X2 U10747 ( .B1(execstage_BusA[4]), .B2(n13164), .A(n5293), .ZN(n5292)
         );
  NOR2_X2 U10748 ( .A1(n3885), .A2(n4037), .ZN(n3884) );
  AOI21_X2 U10749 ( .B1(n13181), .B2(execstage_BusA[15]), .A(n4038), .ZN(n4037) );
  NOR2_X2 U10750 ( .A1(n3560), .A2(n3737), .ZN(n3559) );
  AOI21_X2 U10751 ( .B1(n13181), .B2(execstage_BusA[17]), .A(n3738), .ZN(n3737) );
  NOR2_X2 U10752 ( .A1(n3832), .A2(n3981), .ZN(n3831) );
  AOI21_X2 U10753 ( .B1(execstage_BusA[4]), .B2(n13111), .A(n3982), .ZN(n3981)
         );
  NOR2_X2 U10754 ( .A1(n3676), .A2(n3828), .ZN(n3675) );
  AOI21_X2 U10755 ( .B1(execstage_BusA[4]), .B2(n16431), .A(n3829), .ZN(n3828)
         );
  NOR2_X2 U10756 ( .A1(n3478), .A2(n3672), .ZN(n3477) );
  AOI21_X2 U10757 ( .B1(execstage_BusA[4]), .B2(n16433), .A(n3673), .ZN(n3672)
         );
  NOR2_X2 U10758 ( .A1(n3821), .A2(n16192), .ZN(n3820) );
  OAI21_X2 U10759 ( .B1(n13793), .B2(n3480), .A(n3975), .ZN(n3974) );
  INV_X4 U10760 ( .A(n8693), .ZN(n13119) );
  OAI21_X2 U10761 ( .B1(n8749), .B2(n13763), .A(n312), .ZN(n8302) );
  OAI21_X2 U10762 ( .B1(n8727), .B2(n13763), .A(n312), .ZN(n8304) );
  OAI21_X2 U10763 ( .B1(n8748), .B2(n13763), .A(n312), .ZN(n8306) );
  OAI21_X2 U10764 ( .B1(n13189), .B2(n8731), .A(n3752), .ZN(n3751) );
  OAI21_X2 U10765 ( .B1(n13201), .B2(n8731), .A(n3903), .ZN(n3902) );
  OAI21_X2 U10766 ( .B1(n2869), .B2(n8653), .A(n4196), .ZN(n4195) );
  OAI21_X2 U10767 ( .B1(n2869), .B2(n8733), .A(n3584), .ZN(n3583) );
  INV_X4 U10768 ( .A(n8715), .ZN(n13116) );
  NAND3_X2 U10769 ( .A1(execstage_BusA[21]), .A2(n13191), .A3(n4194), .ZN(
        n4072) );
  INV_X4 U10770 ( .A(n8739), .ZN(n13115) );
  NOR2_X2 U10771 ( .A1(n8717), .A2(n13762), .ZN(n8278) );
  NOR2_X2 U10772 ( .A1(n8726), .A2(n13761), .ZN(n8305) );
  NAND3_X2 U10773 ( .A1(execstage_BusA[8]), .A2(n13176), .A3(n16497), .ZN(
        n5770) );
  NOR2_X2 U10774 ( .A1(n8742), .A2(n13762), .ZN(n8277) );
  NOR2_X2 U10775 ( .A1(n8718), .A2(n13762), .ZN(n8275) );
  NOR2_X2 U10776 ( .A1(n8750), .A2(n13763), .ZN(n8303) );
  NOR2_X2 U10777 ( .A1(n8743), .A2(n13762), .ZN(n8279) );
  NOR2_X2 U10778 ( .A1(n8741), .A2(n13762), .ZN(n8276) );
  NOR2_X2 U10779 ( .A1(n8716), .A2(n13762), .ZN(n8280) );
  NOR2_X2 U10780 ( .A1(n8805), .A2(n13762), .ZN(n8284) );
  NOR2_X2 U10781 ( .A1(n8804), .A2(n13762), .ZN(n8289) );
  NOR2_X2 U10782 ( .A1(n8719), .A2(n13762), .ZN(n8285) );
  NOR2_X2 U10783 ( .A1(n8723), .A2(n13761), .ZN(n8290) );
  NOR2_X2 U10784 ( .A1(n8745), .A2(n13762), .ZN(n8283) );
  NOR2_X2 U10785 ( .A1(n8756), .A2(n13761), .ZN(n8288) );
  NOR2_X2 U10786 ( .A1(n8747), .A2(n13762), .ZN(n8281) );
  NOR2_X2 U10787 ( .A1(n8746), .A2(n13762), .ZN(n8282) );
  NOR2_X2 U10788 ( .A1(n8758), .A2(n13761), .ZN(n8286) );
  NOR2_X2 U10789 ( .A1(n8757), .A2(n13761), .ZN(n8287) );
  NOR2_X2 U10790 ( .A1(n8761), .A2(n13763), .ZN(n8298) );
  NOR2_X2 U10791 ( .A1(n8760), .A2(n13761), .ZN(n8297) );
  NOR2_X2 U10792 ( .A1(n8707), .A2(n13763), .ZN(n8299) );
  NOR2_X2 U10793 ( .A1(n8728), .A2(n13761), .ZN(n8296) );
  NOR2_X2 U10794 ( .A1(n8751), .A2(n13763), .ZN(n8300) );
  NOR2_X2 U10795 ( .A1(n13125), .A2(n8763), .ZN(n8243) );
  NOR2_X2 U10796 ( .A1(n13124), .A2(n8764), .ZN(n8244) );
  NOR2_X2 U10797 ( .A1(n13124), .A2(n8765), .ZN(n8245) );
  NOR2_X2 U10798 ( .A1(n13124), .A2(n8766), .ZN(n8246) );
  NOR2_X2 U10799 ( .A1(n13124), .A2(n8767), .ZN(n8247) );
  NOR2_X2 U10800 ( .A1(n13124), .A2(n8768), .ZN(n8248) );
  NOR2_X2 U10801 ( .A1(n13124), .A2(n8769), .ZN(n8249) );
  NOR2_X2 U10802 ( .A1(n13124), .A2(n8770), .ZN(n8250) );
  NOR2_X2 U10803 ( .A1(n13124), .A2(n8771), .ZN(n8251) );
  NOR2_X2 U10804 ( .A1(n13124), .A2(n8772), .ZN(n8252) );
  NOR2_X2 U10805 ( .A1(n13124), .A2(n8773), .ZN(n8253) );
  NOR2_X2 U10806 ( .A1(n13124), .A2(n8774), .ZN(n8254) );
  NOR2_X2 U10807 ( .A1(n13123), .A2(n8775), .ZN(n8255) );
  NOR2_X2 U10808 ( .A1(n13123), .A2(n8776), .ZN(n8256) );
  NOR2_X2 U10809 ( .A1(n13123), .A2(n8777), .ZN(n8257) );
  NOR2_X2 U10810 ( .A1(n13123), .A2(n8778), .ZN(n8258) );
  NOR2_X2 U10811 ( .A1(n13123), .A2(n8779), .ZN(n8259) );
  NOR2_X2 U10812 ( .A1(n13123), .A2(n8780), .ZN(n8260) );
  NOR2_X2 U10813 ( .A1(n13123), .A2(n8781), .ZN(n8261) );
  NOR2_X2 U10814 ( .A1(n13123), .A2(n8782), .ZN(n8262) );
  NOR2_X2 U10815 ( .A1(n13123), .A2(n8783), .ZN(n8263) );
  NOR2_X2 U10816 ( .A1(n13123), .A2(n8784), .ZN(n8264) );
  NOR2_X2 U10817 ( .A1(n13125), .A2(n8785), .ZN(n8265) );
  NOR2_X2 U10818 ( .A1(n13125), .A2(n8786), .ZN(n8266) );
  NOR2_X2 U10819 ( .A1(n13125), .A2(n8787), .ZN(n8267) );
  NOR2_X2 U10820 ( .A1(n13125), .A2(n8788), .ZN(n8268) );
  NOR2_X2 U10821 ( .A1(n13125), .A2(n8789), .ZN(n8269) );
  NOR2_X2 U10822 ( .A1(n13125), .A2(n8790), .ZN(n8270) );
  NOR2_X2 U10823 ( .A1(n13125), .A2(n8791), .ZN(n8271) );
  NOR2_X2 U10824 ( .A1(n13124), .A2(n8792), .ZN(n8272) );
  NOR2_X2 U10825 ( .A1(n13123), .A2(n8793), .ZN(n8273) );
  NOR2_X2 U10826 ( .A1(n13123), .A2(n8794), .ZN(n8274) );
  INV_X4 U10827 ( .A(execstage_BusA[2]), .ZN(n13793) );
  NOR2_X2 U10828 ( .A1(n4639), .A2(n4753), .ZN(n4638) );
  AOI21_X2 U10829 ( .B1(n13203), .B2(execstage_BusA[18]), .A(n16378), .ZN(
        n4753) );
  INV_X4 U10830 ( .A(n8708), .ZN(n13788) );
  OAI21_X2 U10831 ( .B1(n16393), .B2(n4061), .A(n4062), .ZN(n4059) );
  INV_X4 U10832 ( .A(n8740), .ZN(n13791) );
  AOI222_X1 U10833 ( .A1(n3807), .A2(n2913), .B1(n3808), .B2(n3809), .C1(
        n16427), .C2(n3810), .ZN(n3795) );
  AOI222_X1 U10834 ( .A1(decode_regfile_N136), .A2(n13754), .B1(n13751), .B2(
        n16564), .C1(decode_regfile_N104), .C2(n13748), .ZN(n384) );
  AOI222_X1 U10835 ( .A1(decode_regfile_N135), .A2(n13754), .B1(n13751), .B2(
        n16563), .C1(decode_regfile_N103), .C2(n13748), .ZN(n391) );
  AOI222_X1 U10836 ( .A1(decode_regfile_N134), .A2(n13754), .B1(n13751), .B2(
        n16562), .C1(decode_regfile_N102), .C2(n13748), .ZN(n390) );
  AOI222_X1 U10837 ( .A1(decode_regfile_N29), .A2(n13771), .B1(n13768), .B2(
        n16560), .C1(decode_regfile_N61), .C2(n13765), .ZN(n225) );
  AOI222_X1 U10838 ( .A1(decode_regfile_N30), .A2(n13771), .B1(n13768), .B2(
        n16562), .C1(decode_regfile_N62), .C2(n13765), .ZN(n228) );
  AOI222_X1 U10839 ( .A1(decode_regfile_N28), .A2(n13771), .B1(n13768), .B2(
        n16559), .C1(decode_regfile_N60), .C2(n13765), .ZN(n222) );
  NOR2_X2 U10840 ( .A1(n2909), .A2(n8733), .ZN(n3326) );
  NOR2_X2 U10841 ( .A1(n13148), .A2(n3004), .ZN(n2994) );
  OAI21_X2 U10842 ( .B1(n3000), .B2(n3001), .A(n3002), .ZN(n2996) );
  AOI21_X2 U10843 ( .B1(n3332), .B2(n16481), .A(n16480), .ZN(n3099) );
  NOR2_X2 U10844 ( .A1(n13139), .A2(n5264), .ZN(n5239) );
  INV_X4 U10845 ( .A(n8711), .ZN(n13118) );
  OAI21_X2 U10846 ( .B1(n16372), .B2(n3343), .A(n3344), .ZN(n3072) );
  NOR2_X2 U10847 ( .A1(n8650), .A2(n5264), .ZN(n5616) );
  INV_X4 U10848 ( .A(n8736), .ZN(n13121) );
  INV_X4 U10849 ( .A(n8709), .ZN(n13122) );
  INV_X4 U10850 ( .A(n2869), .ZN(n13202) );
  INV_X4 U10851 ( .A(n3338), .ZN(n13176) );
  INV_X4 U10852 ( .A(n2830), .ZN(n13206) );
  INV_X4 U10853 ( .A(n2869), .ZN(n13203) );
  INV_X4 U10854 ( .A(n8710), .ZN(n13120) );
  INV_X4 U10855 ( .A(n3338), .ZN(n13177) );
  INV_X4 U10856 ( .A(n2869), .ZN(n13204) );
  AOI222_X1 U10857 ( .A1(n16455), .A2(n3237), .B1(n16429), .B2(n3966), .C1(
        n3807), .C2(n3235), .ZN(n3958) );
  AOI222_X1 U10858 ( .A1(n16455), .A2(n3439), .B1(n16435), .B2(n4117), .C1(
        n3807), .C2(n3441), .ZN(n4108) );
  AOI222_X1 U10859 ( .A1(n3807), .A2(n3646), .B1(n16462), .B2(n3806), .C1(
        n16433), .C2(n4263), .ZN(n4255) );
  AOI222_X1 U10860 ( .A1(decode_regfile_N140), .A2(n13753), .B1(n13750), .B2(
        n16568), .C1(decode_regfile_N108), .C2(n13747), .ZN(n370) );
  AOI222_X1 U10861 ( .A1(decode_regfile_N137), .A2(n13754), .B1(n13751), .B2(
        n16565), .C1(decode_regfile_N105), .C2(n13748), .ZN(n385) );
  AOI222_X1 U10862 ( .A1(decode_regfile_N139), .A2(n13754), .B1(n13751), .B2(
        n16567), .C1(decode_regfile_N107), .C2(n13748), .ZN(n387) );
  AOI222_X1 U10863 ( .A1(decode_regfile_N138), .A2(n13754), .B1(n13751), .B2(
        n16566), .C1(decode_regfile_N106), .C2(n13748), .ZN(n386) );
  AOI222_X1 U10864 ( .A1(decode_regfile_N32), .A2(n13771), .B1(n13768), .B2(
        n16564), .C1(decode_regfile_N64), .C2(n13765), .ZN(n234) );
  AOI222_X1 U10865 ( .A1(decode_regfile_N33), .A2(n13771), .B1(n13768), .B2(
        n16565), .C1(decode_regfile_N65), .C2(n13765), .ZN(n237) );
  AOI222_X1 U10866 ( .A1(decode_regfile_N34), .A2(n13771), .B1(n13768), .B2(
        n16566), .C1(decode_regfile_N66), .C2(n13765), .ZN(n240) );
  AOI222_X1 U10867 ( .A1(decode_regfile_N31), .A2(n13771), .B1(n13768), .B2(
        n16563), .C1(decode_regfile_N63), .C2(n13765), .ZN(n231) );
  NOR2_X2 U10868 ( .A1(n8737), .A2(n5264), .ZN(n3238) );
  AOI222_X1 U10869 ( .A1(n8818), .A2(execstage_BusA[23]), .B1(n4532), .B2(
        n13783), .C1(n13131), .C2(n4533), .ZN(n4398) );
  AOI211_X2 U10870 ( .C1(n4264), .C2(n4402), .A(n4403), .B(n16458), .ZN(n4401)
         );
  NOR2_X2 U10871 ( .A1(n4205), .A2(n13194), .ZN(n3638) );
  OAI21_X2 U10872 ( .B1(n13193), .B2(n8653), .A(n4490), .ZN(n4489) );
  OAI21_X2 U10873 ( .B1(n13193), .B2(n8731), .A(n4205), .ZN(n4204) );
  OAI21_X2 U10874 ( .B1(n13193), .B2(n8733), .A(n3641), .ZN(n3906) );
  OAI21_X2 U10875 ( .B1(n3036), .B2(n3037), .A(n3038), .ZN(n3033) );
  OAI21_X2 U10876 ( .B1(n3238), .B2(n3592), .A(n3335), .ZN(n3336) );
  NOR2_X2 U10877 ( .A1(n13194), .A2(n8735), .ZN(n3592) );
  INV_X4 U10878 ( .A(n2804), .ZN(n13210) );
  INV_X4 U10879 ( .A(n2748), .ZN(n13216) );
  INV_X4 U10880 ( .A(execstage_BusA[1]), .ZN(n13149) );
  INV_X4 U10881 ( .A(n2830), .ZN(n13207) );
  INV_X4 U10882 ( .A(n2775), .ZN(n13213) );
  INV_X4 U10883 ( .A(n2804), .ZN(n13211) );
  INV_X4 U10884 ( .A(n2775), .ZN(n13214) );
  INV_X4 U10885 ( .A(n2748), .ZN(n13217) );
  INV_X4 U10886 ( .A(n2830), .ZN(n13208) );
  AOI222_X1 U10887 ( .A1(n3807), .A2(n3965), .B1(n16459), .B2(n2816), .C1(
        n13111), .C2(n4545), .ZN(n4540) );
  AOI222_X1 U10888 ( .A1(decode_regfile_N141), .A2(n13753), .B1(n13750), .B2(
        n16569), .C1(decode_regfile_N109), .C2(n13747), .ZN(n371) );
  AOI222_X1 U10889 ( .A1(decode_regfile_N142), .A2(n13753), .B1(n13750), .B2(
        n16570), .C1(decode_regfile_N110), .C2(n13747), .ZN(n375) );
  AOI222_X1 U10890 ( .A1(decode_regfile_N143), .A2(n13753), .B1(n13750), .B2(
        n16571), .C1(decode_regfile_N111), .C2(n13747), .ZN(n373) );
  AOI222_X1 U10891 ( .A1(decode_regfile_N144), .A2(n13753), .B1(n13750), .B2(
        n16255), .C1(decode_regfile_N112), .C2(n13747), .ZN(n383) );
  AOI222_X1 U10892 ( .A1(decode_regfile_N35), .A2(n13772), .B1(n13769), .B2(
        n16567), .C1(decode_regfile_N67), .C2(n13766), .ZN(n243) );
  AOI222_X1 U10893 ( .A1(decode_regfile_N36), .A2(n13772), .B1(n13769), .B2(
        n16568), .C1(decode_regfile_N68), .C2(n13766), .ZN(n246) );
  AOI222_X1 U10894 ( .A1(decode_regfile_N37), .A2(n13772), .B1(n13769), .B2(
        n16569), .C1(decode_regfile_N69), .C2(n13766), .ZN(n249) );
  AOI222_X1 U10895 ( .A1(decode_regfile_N38), .A2(n13772), .B1(n13769), .B2(
        n16570), .C1(decode_regfile_N70), .C2(n13766), .ZN(n252) );
  AOI222_X1 U10896 ( .A1(n13106), .A2(n3648), .B1(n3807), .B2(n3643), .C1(
        n16455), .C2(n3646), .ZN(n4805) );
  AOI222_X1 U10897 ( .A1(n8818), .A2(execstage_BusA[20]), .B1(n4916), .B2(
        n13782), .C1(n13131), .C2(n4917), .ZN(n4804) );
  AOI222_X1 U10898 ( .A1(n16409), .A2(n4811), .B1(n16468), .B2(n3806), .C1(
        n16440), .C2(n16466), .ZN(n4806) );
  AOI222_X1 U10899 ( .A1(n8818), .A2(execstage_BusA[21]), .B1(n4798), .B2(
        n13782), .C1(n13131), .C2(n4799), .ZN(n4677) );
  AOI211_X2 U10900 ( .C1(n4546), .C2(n4681), .A(n4682), .B(n16458), .ZN(n4680)
         );
  AOI222_X1 U10901 ( .A1(n3806), .A2(n2893), .B1(n4114), .B2(n2892), .C1(
        n13105), .C2(n2913), .ZN(n4950) );
  AOI222_X1 U10902 ( .A1(n8818), .A2(execstage_BusA[19]), .B1(n5057), .B2(
        n13782), .C1(n13131), .C2(n5058), .ZN(n4949) );
  AOI211_X2 U10903 ( .C1(n4815), .C2(n4953), .A(n4954), .B(n16458), .ZN(n4952)
         );
  NOR2_X2 U10904 ( .A1(n8658), .A2(n5264), .ZN(n2921) );
  NOR2_X2 U10905 ( .A1(n3070), .A2(n3071), .ZN(n3069) );
  NOR2_X2 U10906 ( .A1(n13212), .A2(n8731), .ZN(n3075) );
  NOR3_X2 U10907 ( .A1(n3083), .A2(n13189), .A3(n8733), .ZN(n3082) );
  OAI21_X2 U10908 ( .B1(n3063), .B2(n3064), .A(n3065), .ZN(n3058) );
  OAI21_X2 U10909 ( .B1(n3114), .B2(n3115), .A(n3116), .ZN(n3111) );
  NOR2_X2 U10910 ( .A1(n8737), .A2(n13193), .ZN(n3085) );
  NOR2_X2 U10911 ( .A1(n8735), .A2(n13173), .ZN(n3090) );
  INV_X4 U10912 ( .A(n3565), .ZN(n13160) );
  INV_X4 U10913 ( .A(n3130), .ZN(n13181) );
  INV_X4 U10914 ( .A(n3555), .ZN(n13163) );
  INV_X4 U10915 ( .A(n3569), .ZN(n13158) );
  INV_X4 U10916 ( .A(n3130), .ZN(n13182) );
  INV_X4 U10917 ( .A(n3565), .ZN(n13161) );
  INV_X4 U10918 ( .A(n3555), .ZN(n13164) );
  AOI222_X1 U10919 ( .A1(decode_regfile_N41), .A2(n13772), .B1(n13769), .B2(
        n16573), .C1(decode_regfile_N73), .C2(n13766), .ZN(n261) );
  AOI222_X1 U10920 ( .A1(decode_regfile_N39), .A2(n13772), .B1(n13769), .B2(
        n16571), .C1(decode_regfile_N71), .C2(n13766), .ZN(n255) );
  AOI222_X1 U10921 ( .A1(decode_regfile_N40), .A2(n13772), .B1(n13769), .B2(
        n16255), .C1(decode_regfile_N72), .C2(n13766), .ZN(n258) );
  AOI222_X1 U10922 ( .A1(decode_regfile_N42), .A2(n13772), .B1(n13769), .B2(
        n16574), .C1(decode_regfile_N74), .C2(n13766), .ZN(n264) );
  AOI222_X1 U10923 ( .A1(n8818), .A2(execstage_BusA[16]), .B1(n5358), .B2(
        n5359), .C1(n13131), .C2(n5360), .ZN(n5273) );
  AOI222_X1 U10924 ( .A1(n5352), .A2(n13783), .B1(n16455), .B2(n3643), .C1(
        n13105), .C2(n3646), .ZN(n5274) );
  AOI222_X1 U10925 ( .A1(n3807), .A2(n3645), .B1(n4388), .B2(n16459), .C1(
        n13107), .C2(n5278), .ZN(n5275) );
  AOI222_X1 U10926 ( .A1(n3806), .A2(n3419), .B1(n4114), .B2(n3395), .C1(
        n13105), .C2(n3235), .ZN(n5064) );
  AOI222_X1 U10927 ( .A1(n8818), .A2(execstage_BusA[18]), .B1(n5162), .B2(
        n13782), .C1(n13131), .C2(n5163), .ZN(n5063) );
  AOI211_X2 U10928 ( .C1(n4957), .C2(n5067), .A(n5068), .B(n16458), .ZN(n5066)
         );
  AOI222_X1 U10929 ( .A1(n3806), .A2(n4944), .B1(n4114), .B2(n4945), .C1(
        n13106), .C2(n3441), .ZN(n5168) );
  AOI222_X1 U10930 ( .A1(n8818), .A2(execstage_BusA[17]), .B1(n5267), .B2(
        n13782), .C1(n13130), .C2(n5268), .ZN(n5167) );
  AOI211_X2 U10931 ( .C1(n5072), .C2(n5171), .A(n5172), .B(n16458), .ZN(n5170)
         );
  NOR2_X2 U10932 ( .A1(n3099), .A2(n3100), .ZN(n3098) );
  NAND3_X2 U10933 ( .A1(execstage_ALU_ra_row2_31_), .A2(n3101), .A3(n13129), 
        .ZN(n3103) );
  OAI21_X2 U10934 ( .B1(n3060), .B2(n3061), .A(n3062), .ZN(n3059) );
  NOR2_X2 U10935 ( .A1(n8653), .A2(n2748), .ZN(n3050) );
  AOI222_X1 U10936 ( .A1(decode_regfile_N147), .A2(n13753), .B1(n13750), .B2(
        n16575), .C1(decode_regfile_N115), .C2(n13747), .ZN(n377) );
  AOI222_X1 U10937 ( .A1(decode_regfile_N146), .A2(n13753), .B1(n13750), .B2(
        n16574), .C1(decode_regfile_N114), .C2(n13747), .ZN(n379) );
  AOI222_X1 U10938 ( .A1(decode_regfile_N145), .A2(n13753), .B1(n13750), .B2(
        n16573), .C1(decode_regfile_N113), .C2(n13747), .ZN(n381) );
  INV_X4 U10939 ( .A(n3293), .ZN(n13179) );
  INV_X4 U10940 ( .A(n3548), .ZN(n13166) );
  INV_X4 U10941 ( .A(n3543), .ZN(n13168) );
  AOI222_X1 U10942 ( .A1(decode_regfile_N148), .A2(n13752), .B1(n13749), .B2(
        n16576), .C1(decode_regfile_N116), .C2(n13746), .ZN(n343) );
  AOI222_X1 U10943 ( .A1(decode_regfile_N151), .A2(n13752), .B1(n13749), .B2(
        n16579), .C1(decode_regfile_N119), .C2(n13746), .ZN(n333) );
  AOI222_X1 U10944 ( .A1(decode_regfile_N44), .A2(n13770), .B1(n13767), .B2(
        n16576), .C1(decode_regfile_N76), .C2(n13764), .ZN(n63) );
  AOI222_X1 U10945 ( .A1(decode_regfile_N43), .A2(n13770), .B1(n13767), .B2(
        n16575), .C1(decode_regfile_N75), .C2(n13764), .ZN(n57) );
  AOI222_X1 U10946 ( .A1(decode_regfile_N45), .A2(n13770), .B1(n13767), .B2(
        n16577), .C1(decode_regfile_N77), .C2(n13764), .ZN(n66) );
  AOI222_X1 U10947 ( .A1(decode_regfile_N150), .A2(n13752), .B1(n13749), .B2(
        n16578), .C1(decode_regfile_N118), .C2(n13746), .ZN(n339) );
  AOI222_X1 U10948 ( .A1(decode_regfile_N149), .A2(n13752), .B1(n13749), .B2(
        n16577), .C1(decode_regfile_N117), .C2(n13746), .ZN(n341) );
  INV_X4 U10949 ( .A(n13107), .ZN(n13108) );
  INV_X4 U10950 ( .A(n13109), .ZN(n13110) );
  NOR2_X2 U10951 ( .A1(n8716), .A2(n8743), .ZN(n2683) );
  AOI222_X1 U10952 ( .A1(decode_regfile_N152), .A2(n13752), .B1(n13749), .B2(
        n16580), .C1(decode_regfile_N120), .C2(n13746), .ZN(n351) );
  AOI222_X1 U10953 ( .A1(decode_regfile_N154), .A2(n13752), .B1(n13749), .B2(
        n16552), .C1(decode_regfile_N122), .C2(n13746), .ZN(n347) );
  AOI222_X1 U10954 ( .A1(decode_regfile_N153), .A2(n13752), .B1(n13749), .B2(
        n16581), .C1(decode_regfile_N121), .C2(n13746), .ZN(n349) );
  AOI222_X1 U10955 ( .A1(decode_regfile_N46), .A2(n13770), .B1(n13767), .B2(
        n16578), .C1(decode_regfile_N78), .C2(n13764), .ZN(n69) );
  AOI222_X1 U10956 ( .A1(decode_regfile_N48), .A2(n13770), .B1(n13767), .B2(
        n16580), .C1(decode_regfile_N80), .C2(n13764), .ZN(n75) );
  AOI222_X1 U10957 ( .A1(decode_regfile_N47), .A2(n13770), .B1(n13767), .B2(
        n16579), .C1(decode_regfile_N79), .C2(n13764), .ZN(n72) );
  AOI211_X2 U10958 ( .C1(n2683), .C2(n16604), .A(n16594), .B(n16597), .ZN(n143) );
  NOR2_X2 U10959 ( .A1(n16601), .A2(n304), .ZN(n299) );
  NOR2_X2 U10960 ( .A1(n8742), .A2(n8717), .ZN(n2684) );
  NAND3_X2 U10961 ( .A1(n2683), .A2(n8717), .A3(n2681), .ZN(n163) );
  NOR3_X2 U10962 ( .A1(n306), .A2(n2669), .A3(n2687), .ZN(n2660) );
  OAI21_X2 U10963 ( .B1(n2688), .B2(n2689), .A(n301), .ZN(n2687) );
  NOR2_X2 U10964 ( .A1(n2685), .A2(n296), .ZN(n2690) );
  NOR2_X2 U10965 ( .A1(n2691), .A2(n2689), .ZN(n304) );
  AOI211_X2 U10966 ( .C1(n16605), .C2(n296), .A(n145), .B(n16595), .ZN(n294)
         );
  INV_X4 U10967 ( .A(n3500), .ZN(n16406) );
  NAND3_X2 U10968 ( .A1(n2686), .A2(n2684), .A3(n296), .ZN(n2666) );
  NAND3_X2 U10969 ( .A1(n2644), .A2(n302), .A3(n2698), .ZN(n284) );
  AOI21_X2 U10970 ( .B1(n16605), .B2(n2683), .A(n304), .ZN(n2698) );
  INV_X4 U10971 ( .A(n3178), .ZN(n16409) );
  NOR2_X2 U10972 ( .A1(n2926), .A2(n2927), .ZN(n2925) );
  NAND3_X2 U10973 ( .A1(n8741), .A2(n8718), .A3(n2684), .ZN(n2688) );
  AOI222_X1 U10974 ( .A1(decode_regfile_N155), .A2(n13752), .B1(n13749), .B2(
        n16553), .C1(decode_regfile_N123), .C2(n13746), .ZN(n345) );
  INV_X4 U10975 ( .A(n3004), .ZN(n16431) );
  OR2_X2 U10976 ( .A1(n286), .A2(n8719), .ZN(n8810) );
  OR2_X2 U10977 ( .A1(n286), .A2(n8805), .ZN(n8811) );
  INV_X4 U10978 ( .A(n2919), .ZN(n13183) );
  NAND3_X2 U10979 ( .A1(n6039), .A2(n6040), .A3(n6041), .ZN(aluout_0[0]) );
  AOI222_X1 U10980 ( .A1(decode_regfile_N52), .A2(n13770), .B1(n13767), .B2(
        n16554), .C1(decode_regfile_N84), .C2(n13764), .ZN(n87) );
  AOI222_X1 U10981 ( .A1(decode_regfile_N51), .A2(n13770), .B1(n13767), .B2(
        n16553), .C1(decode_regfile_N83), .C2(n13764), .ZN(n84) );
  AOI222_X1 U10982 ( .A1(decode_regfile_N50), .A2(n13770), .B1(n13767), .B2(
        n16552), .C1(decode_regfile_N82), .C2(n13764), .ZN(n81) );
  AOI222_X1 U10983 ( .A1(decode_regfile_N49), .A2(n13770), .B1(n13767), .B2(
        n16581), .C1(decode_regfile_N81), .C2(n13764), .ZN(n78) );
  NOR2_X2 U10984 ( .A1(n286), .A2(n8746), .ZN(decode_rs1_3_) );
  NOR2_X2 U10985 ( .A1(n286), .A2(n8747), .ZN(decode_rs1_4_) );
  AOI222_X1 U10986 ( .A1(decode_regfile_N163), .A2(n13753), .B1(n13750), .B2(
        n16582), .C1(decode_regfile_N131), .C2(n13747), .ZN(n361) );
  AOI222_X1 U10987 ( .A1(decode_regfile_N162), .A2(n13753), .B1(n13750), .B2(
        n16572), .C1(decode_regfile_N130), .C2(n13747), .ZN(n363) );
  AOI222_X1 U10988 ( .A1(decode_regfile_N160), .A2(n13753), .B1(n13750), .B2(
        n16558), .C1(decode_regfile_N128), .C2(n13747), .ZN(n367) );
  AOI222_X1 U10989 ( .A1(decode_regfile_N161), .A2(n13753), .B1(n13750), .B2(
        n16561), .C1(decode_regfile_N129), .C2(n13747), .ZN(n365) );
  AOI222_X1 U10990 ( .A1(decode_regfile_N159), .A2(n13752), .B1(n13749), .B2(
        n16557), .C1(decode_regfile_N127), .C2(n13746), .ZN(n353) );
  AOI222_X1 U10991 ( .A1(decode_regfile_N158), .A2(n13752), .B1(n13749), .B2(
        n16556), .C1(decode_regfile_N126), .C2(n13746), .ZN(n355) );
  AOI222_X1 U10992 ( .A1(decode_regfile_N156), .A2(n13752), .B1(n13749), .B2(
        n16554), .C1(decode_regfile_N124), .C2(n13746), .ZN(n359) );
  AOI222_X1 U10993 ( .A1(decode_regfile_N157), .A2(n13752), .B1(n13749), .B2(
        n16555), .C1(decode_regfile_N125), .C2(n13746), .ZN(n357) );
  AOI222_X1 U10994 ( .A1(decode_regfile_N53), .A2(n13770), .B1(n13767), .B2(
        n16555), .C1(decode_regfile_N85), .C2(n13764), .ZN(n91) );
  AOI222_X1 U10995 ( .A1(decode_regfile_N57), .A2(n13771), .B1(n13768), .B2(
        n16561), .C1(decode_regfile_N89), .C2(n13765), .ZN(n103) );
  AOI222_X1 U10996 ( .A1(decode_regfile_N58), .A2(n13771), .B1(n13768), .B2(
        n16572), .C1(decode_regfile_N90), .C2(n13765), .ZN(n106) );
  AOI222_X1 U10997 ( .A1(decode_regfile_N54), .A2(n13770), .B1(n13767), .B2(
        n16556), .C1(decode_regfile_N86), .C2(n13764), .ZN(n94) );
  AOI222_X1 U10998 ( .A1(decode_regfile_N55), .A2(n13771), .B1(n13768), .B2(
        n16557), .C1(decode_regfile_N87), .C2(n13765), .ZN(n97) );
  AOI222_X1 U10999 ( .A1(decode_regfile_N56), .A2(n13771), .B1(n13768), .B2(
        n16558), .C1(decode_regfile_N88), .C2(n13765), .ZN(n100) );
  INV_X4 U11000 ( .A(n3474), .ZN(n16435) );
  AOI21_X2 U11001 ( .B1(n16411), .B2(n6134), .A(n6135), .ZN(n6133) );
  NOR3_X2 U11002 ( .A1(n16388), .A2(n13113), .A3(n8647), .ZN(n6135) );
  NOR2_X2 U11003 ( .A1(n8651), .A2(n13201), .ZN(n6115) );
  INV_X4 U11004 ( .A(n410), .ZN(n13719) );
  INV_X4 U11005 ( .A(n412), .ZN(n13716) );
  INV_X4 U11006 ( .A(n416), .ZN(n13710) );
  INV_X4 U11007 ( .A(n418), .ZN(n13707) );
  INV_X4 U11008 ( .A(n420), .ZN(n13704) );
  INV_X4 U11009 ( .A(n422), .ZN(n13701) );
  INV_X4 U11010 ( .A(n424), .ZN(n13698) );
  INV_X4 U11011 ( .A(n426), .ZN(n13695) );
  INV_X4 U11012 ( .A(n1565), .ZN(n13393) );
  INV_X4 U11013 ( .A(n1567), .ZN(n13390) );
  INV_X4 U11014 ( .A(n1506), .ZN(n13485) );
  INV_X4 U11015 ( .A(n428), .ZN(n13692) );
  INV_X4 U11016 ( .A(n430), .ZN(n13689) );
  INV_X4 U11017 ( .A(n432), .ZN(n13686) );
  INV_X4 U11018 ( .A(n434), .ZN(n13683) );
  INV_X4 U11019 ( .A(n438), .ZN(n13677) );
  INV_X4 U11020 ( .A(n440), .ZN(n13674) );
  INV_X4 U11021 ( .A(n442), .ZN(n13671) );
  INV_X4 U11022 ( .A(n444), .ZN(n13668) );
  INV_X4 U11023 ( .A(n446), .ZN(n13665) );
  INV_X4 U11024 ( .A(n448), .ZN(n13662) );
  INV_X4 U11025 ( .A(n450), .ZN(n13659) );
  INV_X4 U11026 ( .A(n452), .ZN(n13656) );
  INV_X4 U11027 ( .A(n454), .ZN(n13653) );
  INV_X4 U11028 ( .A(n456), .ZN(n13650) );
  INV_X4 U11029 ( .A(n395), .ZN(n13745) );
  INV_X4 U11030 ( .A(n398), .ZN(n13737) );
  INV_X4 U11031 ( .A(n400), .ZN(n13734) );
  INV_X4 U11032 ( .A(n402), .ZN(n13731) );
  INV_X4 U11033 ( .A(n404), .ZN(n13728) );
  INV_X4 U11034 ( .A(n406), .ZN(n13725) );
  INV_X4 U11035 ( .A(n408), .ZN(n13722) );
  INV_X4 U11036 ( .A(n414), .ZN(n13713) );
  INV_X4 U11037 ( .A(n436), .ZN(n13680) );
  INV_X4 U11038 ( .A(n458), .ZN(n13647) );
  INV_X4 U11039 ( .A(n1521), .ZN(n13459) );
  INV_X4 U11040 ( .A(n1523), .ZN(n13456) );
  INV_X4 U11041 ( .A(n1527), .ZN(n13450) );
  INV_X4 U11042 ( .A(n1529), .ZN(n13447) );
  INV_X4 U11043 ( .A(n1531), .ZN(n13444) );
  INV_X4 U11044 ( .A(n1533), .ZN(n13441) );
  INV_X4 U11045 ( .A(n1535), .ZN(n13438) );
  INV_X4 U11046 ( .A(n1537), .ZN(n13435) );
  INV_X4 U11047 ( .A(n1539), .ZN(n13432) );
  INV_X4 U11048 ( .A(n1541), .ZN(n13429) );
  INV_X4 U11049 ( .A(n1543), .ZN(n13426) );
  INV_X4 U11050 ( .A(n1545), .ZN(n13423) );
  INV_X4 U11051 ( .A(n1549), .ZN(n13417) );
  INV_X4 U11052 ( .A(n1551), .ZN(n13414) );
  INV_X4 U11053 ( .A(n1553), .ZN(n13411) );
  INV_X4 U11054 ( .A(n1555), .ZN(n13408) );
  INV_X4 U11055 ( .A(n1557), .ZN(n13405) );
  INV_X4 U11056 ( .A(n1559), .ZN(n13402) );
  INV_X4 U11057 ( .A(n1561), .ZN(n13399) );
  INV_X4 U11058 ( .A(n1563), .ZN(n13396) );
  INV_X4 U11059 ( .A(n1509), .ZN(n13477) );
  INV_X4 U11060 ( .A(n1511), .ZN(n13474) );
  INV_X4 U11061 ( .A(n1513), .ZN(n13471) );
  INV_X4 U11062 ( .A(n1515), .ZN(n13468) );
  INV_X4 U11063 ( .A(n1517), .ZN(n13465) );
  INV_X4 U11064 ( .A(n1519), .ZN(n13462) );
  INV_X4 U11065 ( .A(n1525), .ZN(n13453) );
  INV_X4 U11066 ( .A(n1547), .ZN(n13420) );
  INV_X4 U11067 ( .A(n1569), .ZN(n13387) );
  NOR2_X2 U11068 ( .A1(execstage_BusA[8]), .A2(n13217), .ZN(n2744) );
  NAND3_X2 U11069 ( .A1(n2684), .A2(n2685), .A3(n2686), .ZN(n280) );
  AOI222_X1 U11070 ( .A1(decode_regfile_N59), .A2(n13771), .B1(n13768), .B2(
        n16582), .C1(decode_regfile_N91), .C2(n13765), .ZN(n109) );
  OAI21_X2 U11071 ( .B1(execstage_BusA[19]), .B2(n3515), .A(n6102), .ZN(n6101)
         );
  NAND3_X2 U11072 ( .A1(n267), .A2(n16174), .A3(n393), .ZN(n8812) );
  NAND3_X2 U11073 ( .A1(n13128), .A2(n16174), .A3(n393), .ZN(n8813) );
  NAND2_X2 U11074 ( .A1(decode_N2), .A2(n393), .ZN(n8814) );
  INV_X4 U11075 ( .A(n3480), .ZN(n16433) );
  NOR2_X2 U11076 ( .A1(n13141), .A2(n3178), .ZN(n3169) );
  INV_X4 U11077 ( .A(decode_rs2_0_), .ZN(n13802) );
  OAI21_X2 U11078 ( .B1(n162), .B2(n8723), .A(n163), .ZN(decode_rs2_0_) );
  OAI21_X2 U11079 ( .B1(n13207), .B2(n13143), .A(n6156), .ZN(n6155) );
  NAND3_X2 U11080 ( .A1(n13189), .A2(n16354), .A3(execstage_BusA[4]), .ZN(
        n6156) );
  NOR2_X2 U11081 ( .A1(n286), .A2(n8745), .ZN(decode_rs1_2_) );
  NOR2_X2 U11082 ( .A1(n3653), .A2(n13192), .ZN(n4114) );
  NOR2_X2 U11083 ( .A1(n3429), .A2(n13190), .ZN(n3808) );
  NAND3_X2 U11084 ( .A1(execstage_ALU_ra_row2_31_), .A2(n13193), .A3(n13129), 
        .ZN(n5811) );
  AOI222_X1 U11085 ( .A1(n4261), .A2(n16471), .B1(n2753), .B2(n8659), .C1(
        n3652), .C2(n8696), .ZN(n2856) );
  NAND3_X2 U11086 ( .A1(n5261), .A2(n5262), .A3(n5263), .ZN(n3441) );
  NAND3_X2 U11087 ( .A1(n5611), .A2(n5054), .A3(n5612), .ZN(n2717) );
  AOI222_X1 U11088 ( .A1(n2907), .A2(n16452), .B1(n13189), .B2(n16385), .C1(
        n2911), .C2(n13191), .ZN(n2906) );
  AOI222_X1 U11089 ( .A1(n2845), .A2(n2846), .B1(n2847), .B2(n16456), .C1(
        n2848), .C2(n2849), .ZN(n2844) );
  NOR2_X2 U11090 ( .A1(n13203), .A2(n2851), .ZN(n2847) );
  OAI21_X2 U11091 ( .B1(n13192), .B2(n13225), .A(n13221), .ZN(n2846) );
  OAI21_X2 U11092 ( .B1(n16451), .B2(n2721), .A(n13219), .ZN(n2848) );
  AOI211_X2 U11093 ( .C1(n3238), .C2(n13193), .A(n3239), .B(n16510), .ZN(n3230) );
  AOI222_X1 U11094 ( .A1(n16469), .A2(n3235), .B1(n16471), .B2(n3236), .C1(
        n8696), .C2(n3237), .ZN(n3232) );
  NOR3_X2 U11095 ( .A1(n3637), .A2(n3638), .A3(n16511), .ZN(n3636) );
  AOI222_X1 U11096 ( .A1(n8659), .A2(n3643), .B1(n13202), .B2(n16474), .C1(
        n16471), .C2(n3645), .ZN(n3635) );
  AOI222_X1 U11097 ( .A1(n16469), .A2(n3646), .B1(n16471), .B2(n3647), .C1(
        n8696), .C2(n3648), .ZN(n3634) );
  AOI222_X1 U11098 ( .A1(n13191), .A2(n3430), .B1(n16383), .B2(n13189), .C1(
        n16452), .C2(n3432), .ZN(n3428) );
  NOR2_X2 U11099 ( .A1(n4394), .A2(n4248), .ZN(n6161) );
  NOR2_X2 U11100 ( .A1(n3231), .A2(n3653), .ZN(n3220) );
  OAI21_X2 U11101 ( .B1(n8744), .B2(n13184), .A(n5608), .ZN(n3445) );
  NAND3_X2 U11102 ( .A1(execstage_ALU_ra_row2_31_), .A2(n13103), .A3(n3806), 
        .ZN(n3955) );
  OAI21_X2 U11103 ( .B1(n13171), .B2(n8744), .A(n3243), .ZN(n3245) );
  OAI21_X2 U11104 ( .B1(n13197), .B2(n5619), .A(n4933), .ZN(n4941) );
  OAI21_X2 U11105 ( .B1(n16323), .B2(n2721), .A(n13219), .ZN(n2713) );
  OAI21_X2 U11106 ( .B1(n8744), .B2(n13194), .A(n5608), .ZN(n3443) );
  NOR2_X2 U11107 ( .A1(n8738), .A2(n3209), .ZN(n3207) );
  NAND3_X2 U11108 ( .A1(n4100), .A2(n3241), .A3(n6015), .ZN(n4667) );
  OAI21_X2 U11109 ( .B1(n3244), .B2(n3220), .A(n3652), .ZN(n3651) );
  AOI21_X2 U11110 ( .B1(n16534), .B2(n13194), .A(n3638), .ZN(n6017) );
  AOI21_X2 U11111 ( .B1(n16535), .B2(n13194), .A(n16505), .ZN(n6176) );
  NAND3_X2 U11112 ( .A1(n4389), .A2(n3640), .A3(n6180), .ZN(n4261) );
  AOI21_X2 U11113 ( .B1(n16538), .B2(n13194), .A(n16508), .ZN(n6180) );
  OAI21_X2 U11114 ( .B1(n13193), .B2(n2880), .A(n4933), .ZN(n4932) );
  OAI21_X2 U11115 ( .B1(n13193), .B2(n3408), .A(n3409), .ZN(n3407) );
  OAI21_X2 U11116 ( .B1(n8658), .B2(n13219), .A(n16444), .ZN(n3228) );
  OAI21_X2 U11117 ( .B1(n8735), .B2(n13219), .A(n16444), .ZN(n3633) );
  NOR2_X2 U11118 ( .A1(n13793), .A2(n2970), .ZN(n2968) );
  NAND4_X2 U11119 ( .A1(n266), .A2(n267), .A3(n16175), .A4(n16547), .ZN(n8815)
         );
  NAND4_X2 U11120 ( .A1(n13128), .A2(n266), .A3(n16175), .A4(n16547), .ZN(
        n8816) );
  NAND3_X2 U11121 ( .A1(n266), .A2(n16547), .A3(decode_N4), .ZN(n8817) );
  INV_X4 U11122 ( .A(n8818), .ZN(n13219) );
  INV_X4 U11123 ( .A(n8818), .ZN(n13220) );
  NAND2_X2 U11124 ( .A1(n6045), .A2(n8720), .ZN(n2896) );
  INV_X4 U11125 ( .A(n13784), .ZN(n13782) );
  INV_X4 U11126 ( .A(execstage_ALU_N160), .ZN(n13784) );
  INV_X4 U11127 ( .A(n13784), .ZN(n13783) );
  INV_X4 U11128 ( .A(rgwrite_jalout), .ZN(n13781) );
  NOR2_X2 U11129 ( .A1(n3222), .A2(n13192), .ZN(n3806) );
  INV_X4 U11130 ( .A(decode_rs2_1_), .ZN(n13800) );
  OAI21_X2 U11131 ( .B1(n162), .B2(n8804), .A(n163), .ZN(decode_rs2_1_) );
  OAI21_X2 U11132 ( .B1(n162), .B2(n8757), .A(n163), .ZN(decode_rs2_3_) );
  OAI21_X2 U11133 ( .B1(n162), .B2(n8758), .A(n163), .ZN(decode_rs2_4_) );
  INV_X4 U11134 ( .A(decode_rs2_2_), .ZN(n13799) );
  OAI21_X2 U11135 ( .B1(n162), .B2(n8756), .A(n163), .ZN(decode_rs2_2_) );
  NOR3_X2 U11136 ( .A1(n19), .A2(n159), .A3(n160), .ZN(execstage_register_N50)
         );
  NOR2_X2 U11137 ( .A1(n2909), .A2(n3222), .ZN(n2733) );
  INV_X4 U11138 ( .A(n8722), .ZN(n13114) );
  NOR2_X2 U11139 ( .A1(n149), .A2(n137), .ZN(n138) );
  NOR2_X2 U11140 ( .A1(n8729), .A2(n8752), .ZN(n836) );
  NAND3_X2 U11141 ( .A1(n2679), .A2(n8743), .A3(n2697), .ZN(n149) );
  NOR2_X2 U11142 ( .A1(n8748), .A2(n8726), .ZN(n2658) );
  NAND3_X2 U11143 ( .A1(n2697), .A2(n2679), .A3(n2683), .ZN(n220) );
  NOR2_X2 U11144 ( .A1(n2657), .A2(n2658), .ZN(n2646) );
  NOR2_X2 U11145 ( .A1(n2373), .A2(n8753), .ZN(n1939) );
  NOR2_X2 U11146 ( .A1(n8753), .A2(n1270), .ZN(n835) );
  NOR3_X2 U11147 ( .A1(n202), .A2(n191), .A3(n20), .ZN(execstage_register_N13)
         );
  NAND3_X2 U11148 ( .A1(n2697), .A2(n2679), .A3(n16599), .ZN(n2700) );
  NOR2_X2 U11149 ( .A1(n13805), .A2(n8717), .ZN(execstage_register_N180) );
  NOR2_X2 U11150 ( .A1(n13806), .A2(n8726), .ZN(execstage_register_N20) );
  NOR2_X2 U11151 ( .A1(n13806), .A2(n8742), .ZN(execstage_register_N181) );
  NOR2_X2 U11152 ( .A1(n13806), .A2(n8727), .ZN(execstage_register_N21) );
  NOR2_X2 U11153 ( .A1(n13806), .A2(n8718), .ZN(execstage_register_N183) );
  NOR2_X2 U11154 ( .A1(n13806), .A2(n8750), .ZN(execstage_register_N22) );
  NOR2_X2 U11155 ( .A1(n13805), .A2(n8743), .ZN(execstage_register_N179) );
  NOR2_X2 U11156 ( .A1(n13806), .A2(n8748), .ZN(execstage_register_N19) );
  NOR2_X2 U11157 ( .A1(n13806), .A2(n8741), .ZN(execstage_register_N182) );
  NOR2_X2 U11158 ( .A1(n13805), .A2(n8716), .ZN(execstage_register_N178) );
  NOR2_X2 U11159 ( .A1(n13806), .A2(n8749), .ZN(execstage_register_N23) );
  NOR2_X2 U11160 ( .A1(n13807), .A2(n161), .ZN(execstage_register_N5) );
  NOR2_X2 U11161 ( .A1(n13806), .A2(n8761), .ZN(execstage_register_N27) );
  NOR2_X2 U11162 ( .A1(n13806), .A2(n8760), .ZN(execstage_register_N28) );
  NOR2_X2 U11163 ( .A1(n13806), .A2(n8707), .ZN(execstage_register_N26) );
  NOR2_X2 U11164 ( .A1(n13806), .A2(n8751), .ZN(execstage_register_N25) );
  NOR2_X2 U11165 ( .A1(n13806), .A2(n8728), .ZN(execstage_register_N29) );
  NOR2_X2 U11166 ( .A1(n13805), .A2(n8763), .ZN(execstage_register_N151) );
  NOR2_X2 U11167 ( .A1(n13805), .A2(n8764), .ZN(execstage_register_N150) );
  NOR2_X2 U11168 ( .A1(n13805), .A2(n8765), .ZN(execstage_register_N149) );
  NOR2_X2 U11169 ( .A1(n13805), .A2(n8766), .ZN(execstage_register_N148) );
  NOR2_X2 U11170 ( .A1(n13805), .A2(n8767), .ZN(execstage_register_N147) );
  NOR2_X2 U11171 ( .A1(n13805), .A2(n8768), .ZN(execstage_register_N146) );
  NOR2_X2 U11172 ( .A1(n13805), .A2(n8769), .ZN(execstage_register_N145) );
  NOR2_X2 U11173 ( .A1(n13805), .A2(n8770), .ZN(execstage_register_N144) );
  NOR2_X2 U11174 ( .A1(n13805), .A2(n8771), .ZN(execstage_register_N143) );
  NOR2_X2 U11175 ( .A1(stall), .A2(n8772), .ZN(execstage_register_N142) );
  NOR2_X2 U11176 ( .A1(stall), .A2(n8773), .ZN(execstage_register_N141) );
  NOR2_X2 U11177 ( .A1(stall), .A2(n8774), .ZN(execstage_register_N140) );
  NOR2_X2 U11178 ( .A1(stall), .A2(n8775), .ZN(execstage_register_N139) );
  NOR2_X2 U11179 ( .A1(stall), .A2(n8776), .ZN(execstage_register_N138) );
  NOR2_X2 U11180 ( .A1(stall), .A2(n8777), .ZN(execstage_register_N137) );
  NOR2_X2 U11181 ( .A1(stall), .A2(n8778), .ZN(execstage_register_N136) );
  NOR2_X2 U11182 ( .A1(stall), .A2(n8779), .ZN(execstage_register_N135) );
  NOR2_X2 U11183 ( .A1(n13805), .A2(n8780), .ZN(execstage_register_N134) );
  NOR2_X2 U11184 ( .A1(stall), .A2(n8781), .ZN(execstage_register_N133) );
  NOR2_X2 U11185 ( .A1(n13808), .A2(n8782), .ZN(execstage_register_N132) );
  NOR2_X2 U11186 ( .A1(stall), .A2(n8783), .ZN(execstage_register_N131) );
  NOR2_X2 U11187 ( .A1(n13808), .A2(n8784), .ZN(execstage_register_N130) );
  NOR2_X2 U11188 ( .A1(n13804), .A2(n8785), .ZN(execstage_register_N129) );
  NOR2_X2 U11189 ( .A1(stall), .A2(n8786), .ZN(execstage_register_N128) );
  NOR2_X2 U11190 ( .A1(n13804), .A2(n8787), .ZN(execstage_register_N127) );
  NOR2_X2 U11191 ( .A1(n13804), .A2(n8788), .ZN(execstage_register_N126) );
  NOR2_X2 U11192 ( .A1(n13804), .A2(n8789), .ZN(execstage_register_N125) );
  NOR2_X2 U11193 ( .A1(n13804), .A2(n8790), .ZN(execstage_register_N124) );
  NOR2_X2 U11194 ( .A1(n13804), .A2(n8791), .ZN(execstage_register_N123) );
  NOR2_X2 U11195 ( .A1(n13804), .A2(n8792), .ZN(execstage_register_N122) );
  NOR2_X2 U11196 ( .A1(n13804), .A2(n8793), .ZN(execstage_register_N121) );
  NOR2_X2 U11197 ( .A1(n13804), .A2(n8794), .ZN(execstage_register_N120) );
  INV_X4 U11198 ( .A(n8819), .ZN(n13228) );
  INV_X4 U11199 ( .A(n8820), .ZN(n13486) );
  INV_X4 U11200 ( .A(n8821), .ZN(n13488) );
  INV_X4 U11201 ( .A(n8819), .ZN(n13229) );
  INV_X4 U11202 ( .A(n8820), .ZN(n13487) );
  INV_X4 U11203 ( .A(n8821), .ZN(n13489) );
  INV_X4 U11204 ( .A(mem_memtoreg_out), .ZN(n13127) );
  INV_X4 U11205 ( .A(mem_memtoreg_out), .ZN(n13126) );
  AOI211_X2 U11206 ( .C1(n138), .C2(n2651), .A(n284), .B(n16592), .ZN(n2650)
         );
  NAND3_X2 U11207 ( .A1(n2652), .A2(n2648), .A3(n16583), .ZN(n2651) );
  AOI211_X2 U11208 ( .C1(n138), .C2(n2668), .A(n2669), .B(n16589), .ZN(n2667)
         );
  OAI21_X2 U11209 ( .B1(n147), .B2(n2675), .A(n2647), .ZN(n2665) );
  OAI21_X2 U11210 ( .B1(n2659), .B2(n16588), .A(n2660), .ZN(
        decode_decoder_N277) );
  AOI211_X2 U11211 ( .C1(n2658), .C2(n2656), .A(n16585), .B(n2662), .ZN(n2659)
         );
  NAND3_X2 U11212 ( .A1(n8727), .A2(n8750), .A3(n16587), .ZN(n2655) );
  INV_X4 U11213 ( .A(n8822), .ZN(n13756) );
  INV_X4 U11214 ( .A(execstage_ALU_sel), .ZN(n13132) );
  INV_X4 U11215 ( .A(execstage_ALU_sel), .ZN(n13133) );
  INV_X4 U11216 ( .A(n8822), .ZN(n13755) );
  INV_X4 U11217 ( .A(n8823), .ZN(n13776) );
  INV_X4 U11218 ( .A(n8823), .ZN(n13777) );
  INV_X4 U11219 ( .A(n8824), .ZN(n13759) );
  INV_X4 U11220 ( .A(n8824), .ZN(n13758) );
  INV_X4 U11221 ( .A(n8823), .ZN(n13778) );
  INV_X4 U11222 ( .A(n8824), .ZN(n13760) );
  INV_X4 U11223 ( .A(n8822), .ZN(n13757) );
  INV_X4 U11224 ( .A(n8825), .ZN(n13774) );
  INV_X4 U11225 ( .A(n8825), .ZN(n13773) );
  INV_X4 U11226 ( .A(n8825), .ZN(n13775) );
  INV_X4 U11227 ( .A(execstage_ALU_sel), .ZN(n13134) );
  NAND3_X2 U11228 ( .A1(execstage_BusA[25]), .A2(n13191), .A3(n3582), .ZN(
        n3344) );
  NAND3_X2 U11229 ( .A1(n13176), .A2(execstage_BusA[1]), .A3(n5990), .ZN(n5988) );
  NOR2_X2 U11230 ( .A1(n3774), .A2(n3898), .ZN(n3773) );
  AOI21_X2 U11231 ( .B1(n13206), .B2(execstage_BusA[22]), .A(n3899), .ZN(n3898) );
  INV_X4 U11232 ( .A(n2881), .ZN(n13200) );
  NOR2_X2 U11233 ( .A1(n8759), .A2(n13763), .ZN(n8301) );
  NOR2_X2 U11234 ( .A1(n8798), .A2(n13761), .ZN(n8291) );
  NOR2_X2 U11235 ( .A1(n8799), .A2(n13761), .ZN(n8292) );
  NOR2_X2 U11236 ( .A1(n8800), .A2(n13761), .ZN(n8293) );
  NOR2_X2 U11237 ( .A1(n8801), .A2(n13761), .ZN(n8294) );
  NOR2_X2 U11238 ( .A1(n8802), .A2(n13761), .ZN(n8295) );
  INV_X4 U11239 ( .A(n5264), .ZN(n13102) );
  OAI22_X2 U11240 ( .A1(execstage_Imm32[0]), .A2(n13787), .B1(n13788), .B2(
        busB_1[0]), .ZN(n5264) );
  NOR2_X2 U11241 ( .A1(n3913), .A2(n4055), .ZN(n3912) );
  AOI21_X2 U11242 ( .B1(n13177), .B2(execstage_BusA[24]), .A(n16391), .ZN(
        n4055) );
  AOI222_X1 U11243 ( .A1(n3945), .A2(n13783), .B1(n16455), .B2(n2916), .C1(
        n13106), .C2(n2915), .ZN(n3794) );
  AOI211_X2 U11244 ( .C1(n3659), .C2(n3797), .A(n16445), .B(n3799), .ZN(n3796)
         );
  INV_X4 U11245 ( .A(n2909), .ZN(n13188) );
  NAND3_X2 U11246 ( .A1(n3422), .A2(n3423), .A3(n3424), .ZN(aluout_0[29]) );
  AOI211_X2 U11247 ( .C1(n13218), .C2(execstage_BusA[29]), .A(n3425), .B(n3426), .ZN(n3424) );
  AOI222_X1 U11248 ( .A1(n3244), .A2(n3443), .B1(n3390), .B2(n3444), .C1(n3220), .C2(n3445), .ZN(n3423) );
  INV_X4 U11249 ( .A(execstage_BusA[20]), .ZN(n13117) );
  INV_X4 U11250 ( .A(n3569), .ZN(n13156) );
  AOI222_X1 U11251 ( .A1(n8818), .A2(execstage_BusA[26]), .B1(n3808), .B2(
        n4104), .C1(n13131), .C2(n4105), .ZN(n3956) );
  AOI222_X1 U11252 ( .A1(n3806), .A2(n16461), .B1(n13106), .B2(n3236), .C1(
        n4096), .C2(n13783), .ZN(n3957) );
  AOI211_X2 U11253 ( .C1(n3811), .C2(n3960), .A(n3961), .B(n16458), .ZN(n3959)
         );
  AOI222_X1 U11254 ( .A1(n3806), .A2(n2734), .B1(n3808), .B2(n2732), .C1(
        n13105), .C2(n3440), .ZN(n4107) );
  AOI222_X1 U11255 ( .A1(n13218), .A2(execstage_BusA[25]), .B1(n4247), .B2(
        n13783), .C1(n13131), .C2(n4248), .ZN(n4106) );
  AOI211_X2 U11256 ( .C1(n3967), .C2(n4110), .A(n4111), .B(n16458), .ZN(n4109)
         );
  AOI222_X1 U11257 ( .A1(n13105), .A2(n3647), .B1(n16455), .B2(n3648), .C1(
        n3808), .C2(n16465), .ZN(n4254) );
  AOI222_X1 U11258 ( .A1(n8818), .A2(execstage_BusA[24]), .B1(n4393), .B2(
        n13782), .C1(n13131), .C2(n4394), .ZN(n4253) );
  AOI211_X2 U11259 ( .C1(n4118), .C2(n4257), .A(n4258), .B(n16458), .ZN(n4256)
         );
  NAND3_X2 U11260 ( .A1(n3238), .A2(n13197), .A3(execstage_BusA[28]), .ZN(
        n3335) );
  AOI222_X1 U11261 ( .A1(n8818), .A2(execstage_BusA[22]), .B1(n4672), .B2(
        n13782), .C1(n13131), .C2(n4673), .ZN(n4538) );
  AOI211_X2 U11262 ( .C1(n4408), .C2(n4542), .A(n4543), .B(n16458), .ZN(n4541)
         );
  INV_X4 U11263 ( .A(n3145), .ZN(n13107) );
  OAI22_X2 U11264 ( .A1(execstage_Imm32[16]), .A2(n13786), .B1(n13788), .B2(
        busB_1[16]), .ZN(n3145) );
  INV_X4 U11265 ( .A(n3529), .ZN(n13113) );
  OAI22_X2 U11266 ( .A1(execstage_Imm32[17]), .A2(n13785), .B1(
        execstage_ALUSrc), .B2(busB_1[17]), .ZN(n3529) );
  INV_X4 U11267 ( .A(n3201), .ZN(n13109) );
  OAI22_X2 U11268 ( .A1(execstage_Imm32[18]), .A2(n13785), .B1(n13788), .B2(
        busB_1[18]), .ZN(n3201) );
  INV_X4 U11269 ( .A(n3515), .ZN(n13112) );
  OAI22_X2 U11270 ( .A1(execstage_Imm32[19]), .A2(n13785), .B1(
        execstage_ALUSrc), .B2(busB_1[19]), .ZN(n3515) );
  OAI22_X2 U11271 ( .A1(execstage_Imm32[21]), .A2(n13785), .B1(
        execstage_ALUSrc), .B2(busB_1[21]), .ZN(n3500) );
  NOR2_X2 U11272 ( .A1(instruction_1[27]), .A2(instruction_1[26]), .ZN(n296)
         );
  NOR2_X2 U11273 ( .A1(instruction_1[30]), .A2(instruction_1[28]), .ZN(n2697)
         );
  NOR2_X2 U11274 ( .A1(instruction_1[31]), .A2(instruction_1[29]), .ZN(n2679)
         );
  NOR2_X2 U11275 ( .A1(n8741), .A2(instruction_1[31]), .ZN(n2686) );
  NOR2_X2 U11276 ( .A1(n8716), .A2(instruction_1[27]), .ZN(n2685) );
  OAI21_X2 U11277 ( .B1(n2696), .B2(n16595), .A(n8742), .ZN(n161) );
  NOR3_X2 U11278 ( .A1(n8718), .A2(instruction_1[30]), .A3(n2690), .ZN(n2696)
         );
  NAND3_X2 U11279 ( .A1(instruction_1[28]), .A2(n16599), .A3(n2681), .ZN(n302)
         );
  NAND3_X2 U11280 ( .A1(n2681), .A2(instruction_1[28]), .A3(n296), .ZN(n2644)
         );
  NAND3_X2 U11281 ( .A1(instruction_1[28]), .A2(n2683), .A3(n2681), .ZN(n2649)
         );
  NAND3_X2 U11282 ( .A1(n2697), .A2(n8718), .A3(instruction_1[29]), .ZN(n2691)
         );
  NAND3_X2 U11283 ( .A1(instruction_1[29]), .A2(n8717), .A3(n2686), .ZN(n2695)
         );
  OAI22_X2 U11284 ( .A1(execstage_Imm32[20]), .A2(n13785), .B1(n13788), .B2(
        busB_1[20]), .ZN(n3178) );
  OAI22_X2 U11285 ( .A1(execstage_Imm32[23]), .A2(n13787), .B1(n13788), .B2(
        busB_1[23]), .ZN(n3004) );
  INV_X4 U11286 ( .A(n3494), .ZN(n13111) );
  OAI22_X2 U11287 ( .A1(execstage_Imm32[22]), .A2(n13785), .B1(n13788), .B2(
        busB_1[22]), .ZN(n3494) );
  OAI22_X2 U11288 ( .A1(execstage_Imm32[26]), .A2(n13786), .B1(n13788), .B2(
        busB_1[26]), .ZN(n2946) );
  AOI222_X1 U11289 ( .A1(execstage_BusA[30]), .A2(n6128), .B1(n16436), .B2(
        n6129), .C1(n16422), .C2(n6131), .ZN(n6127) );
  AOI21_X2 U11290 ( .B1(n6085), .B2(n6086), .A(n6087), .ZN(n6084) );
  AOI21_X2 U11291 ( .B1(n6058), .B2(n6059), .A(execstage_AluCtrl[2]), .ZN(
        n6053) );
  NOR2_X2 U11292 ( .A1(execstage_AluCtrl[1]), .A2(n6057), .ZN(n6058) );
  AOI21_X2 U11293 ( .B1(execstage_AluCtrl[1]), .B2(n6060), .A(n8660), .ZN(
        n6052) );
  OAI21_X2 U11294 ( .B1(execstage_AluCtrl[0]), .B2(n6059), .A(n6061), .ZN(
        n6060) );
  NAND3_X2 U11295 ( .A1(n6062), .A2(n6056), .A3(execstage_AluCtrl[0]), .ZN(
        n6061) );
  NOR3_X2 U11296 ( .A1(n13193), .A2(execstage_BusA[1]), .A3(n3418), .ZN(n6125)
         );
  OAI21_X2 U11297 ( .B1(n13718), .B2(n13545), .A(n1111), .ZN(n6227) );
  OAI21_X2 U11298 ( .B1(n13715), .B2(n13546), .A(n1112), .ZN(n6228) );
  OAI21_X2 U11299 ( .B1(n13709), .B2(n13546), .A(n1114), .ZN(n6229) );
  OAI21_X2 U11300 ( .B1(n13706), .B2(n13546), .A(n1115), .ZN(n6230) );
  OAI21_X2 U11301 ( .B1(n13703), .B2(n13546), .A(n1116), .ZN(n6231) );
  OAI21_X2 U11302 ( .B1(n13700), .B2(n13546), .A(n1117), .ZN(n6232) );
  OAI21_X2 U11303 ( .B1(n13697), .B2(n13546), .A(n1118), .ZN(n6233) );
  OAI21_X2 U11304 ( .B1(n13694), .B2(n13546), .A(n1119), .ZN(n6234) );
  OAI21_X2 U11305 ( .B1(n13691), .B2(n13547), .A(n1120), .ZN(n6235) );
  OAI21_X2 U11306 ( .B1(n13688), .B2(n13547), .A(n1121), .ZN(n6236) );
  OAI21_X2 U11307 ( .B1(n13685), .B2(n13546), .A(n1122), .ZN(n6237) );
  OAI21_X2 U11308 ( .B1(n13682), .B2(n13547), .A(n1123), .ZN(n6238) );
  OAI21_X2 U11309 ( .B1(n13676), .B2(n13547), .A(n1125), .ZN(n6239) );
  OAI21_X2 U11310 ( .B1(n13673), .B2(n13547), .A(n1126), .ZN(n6240) );
  OAI21_X2 U11311 ( .B1(n13670), .B2(n13547), .A(n1127), .ZN(n6241) );
  OAI21_X2 U11312 ( .B1(n13667), .B2(n13547), .A(n1128), .ZN(n6242) );
  OAI21_X2 U11313 ( .B1(n13664), .B2(n13546), .A(n1129), .ZN(n6243) );
  OAI21_X2 U11314 ( .B1(n13661), .B2(n13546), .A(n1130), .ZN(n6244) );
  OAI21_X2 U11315 ( .B1(n13658), .B2(n13546), .A(n1131), .ZN(n6245) );
  OAI21_X2 U11316 ( .B1(n13655), .B2(n13545), .A(n1132), .ZN(n6246) );
  OAI21_X2 U11317 ( .B1(n13652), .B2(n13545), .A(n1133), .ZN(n6247) );
  OAI21_X2 U11318 ( .B1(n13649), .B2(n13545), .A(n1134), .ZN(n6248) );
  OAI21_X2 U11319 ( .B1(n13744), .B2(n13545), .A(n1104), .ZN(n6249) );
  OAI21_X2 U11320 ( .B1(n13736), .B2(n13545), .A(n1105), .ZN(n6250) );
  OAI21_X2 U11321 ( .B1(n13733), .B2(n13545), .A(n1106), .ZN(n6251) );
  OAI21_X2 U11322 ( .B1(n13730), .B2(n13545), .A(n1107), .ZN(n6252) );
  OAI21_X2 U11323 ( .B1(n13727), .B2(n13545), .A(n1108), .ZN(n6253) );
  OAI21_X2 U11324 ( .B1(n13724), .B2(n13545), .A(n1109), .ZN(n6254) );
  OAI21_X2 U11325 ( .B1(n13721), .B2(n13545), .A(n1110), .ZN(n6255) );
  OAI21_X2 U11326 ( .B1(n13712), .B2(n13546), .A(n1113), .ZN(n6256) );
  OAI21_X2 U11327 ( .B1(n13679), .B2(n13547), .A(n1124), .ZN(n6257) );
  OAI21_X2 U11328 ( .B1(n13646), .B2(n13545), .A(n1135), .ZN(n6258) );
  OAI21_X2 U11329 ( .B1(n13717), .B2(n13615), .A(n639), .ZN(n6291) );
  OAI21_X2 U11330 ( .B1(n13714), .B2(n13616), .A(n640), .ZN(n6292) );
  OAI21_X2 U11331 ( .B1(n13708), .B2(n13616), .A(n642), .ZN(n6293) );
  OAI21_X2 U11332 ( .B1(n13705), .B2(n13616), .A(n643), .ZN(n6294) );
  OAI21_X2 U11333 ( .B1(n13702), .B2(n13616), .A(n644), .ZN(n6295) );
  OAI21_X2 U11334 ( .B1(n13699), .B2(n13616), .A(n645), .ZN(n6296) );
  OAI21_X2 U11335 ( .B1(n13696), .B2(n13616), .A(n646), .ZN(n6297) );
  OAI21_X2 U11336 ( .B1(n13693), .B2(n13616), .A(n647), .ZN(n6298) );
  OAI21_X2 U11337 ( .B1(n13690), .B2(n13617), .A(n648), .ZN(n6299) );
  OAI21_X2 U11338 ( .B1(n13687), .B2(n13617), .A(n649), .ZN(n6300) );
  OAI21_X2 U11339 ( .B1(n13684), .B2(n13616), .A(n650), .ZN(n6301) );
  OAI21_X2 U11340 ( .B1(n13681), .B2(n13617), .A(n651), .ZN(n6302) );
  OAI21_X2 U11341 ( .B1(n13675), .B2(n13617), .A(n653), .ZN(n6303) );
  OAI21_X2 U11342 ( .B1(n13672), .B2(n13617), .A(n654), .ZN(n6304) );
  OAI21_X2 U11343 ( .B1(n13669), .B2(n13617), .A(n655), .ZN(n6305) );
  OAI21_X2 U11344 ( .B1(n13666), .B2(n13617), .A(n656), .ZN(n6306) );
  OAI21_X2 U11345 ( .B1(n13663), .B2(n13616), .A(n657), .ZN(n6307) );
  OAI21_X2 U11346 ( .B1(n13660), .B2(n13616), .A(n658), .ZN(n6308) );
  OAI21_X2 U11347 ( .B1(n13657), .B2(n13616), .A(n659), .ZN(n6309) );
  OAI21_X2 U11348 ( .B1(n13654), .B2(n13615), .A(n660), .ZN(n6310) );
  OAI21_X2 U11349 ( .B1(n13651), .B2(n13615), .A(n661), .ZN(n6311) );
  OAI21_X2 U11350 ( .B1(n13648), .B2(n13615), .A(n662), .ZN(n6312) );
  OAI21_X2 U11351 ( .B1(n13743), .B2(n13615), .A(n632), .ZN(n6313) );
  OAI21_X2 U11352 ( .B1(n13735), .B2(n13615), .A(n633), .ZN(n6314) );
  OAI21_X2 U11353 ( .B1(n13732), .B2(n13615), .A(n634), .ZN(n6315) );
  OAI21_X2 U11354 ( .B1(n13729), .B2(n13615), .A(n635), .ZN(n6316) );
  OAI21_X2 U11355 ( .B1(n13726), .B2(n13615), .A(n636), .ZN(n6317) );
  OAI21_X2 U11356 ( .B1(n13723), .B2(n13615), .A(n637), .ZN(n6318) );
  OAI21_X2 U11357 ( .B1(n13720), .B2(n13615), .A(n638), .ZN(n6319) );
  OAI21_X2 U11358 ( .B1(n13711), .B2(n13616), .A(n641), .ZN(n6320) );
  OAI21_X2 U11359 ( .B1(n13678), .B2(n13617), .A(n652), .ZN(n6321) );
  OAI21_X2 U11360 ( .B1(n13645), .B2(n13615), .A(n663), .ZN(n6322) );
  OAI21_X2 U11361 ( .B1(n13717), .B2(n13625), .A(n573), .ZN(n6355) );
  OAI21_X2 U11362 ( .B1(n13714), .B2(n13626), .A(n574), .ZN(n6356) );
  OAI21_X2 U11363 ( .B1(n13708), .B2(n13626), .A(n576), .ZN(n6357) );
  OAI21_X2 U11364 ( .B1(n13705), .B2(n13626), .A(n577), .ZN(n6358) );
  OAI21_X2 U11365 ( .B1(n13702), .B2(n13626), .A(n578), .ZN(n6359) );
  OAI21_X2 U11366 ( .B1(n13699), .B2(n13626), .A(n579), .ZN(n6360) );
  OAI21_X2 U11367 ( .B1(n13696), .B2(n13626), .A(n580), .ZN(n6361) );
  OAI21_X2 U11368 ( .B1(n13693), .B2(n13626), .A(n581), .ZN(n6362) );
  OAI21_X2 U11369 ( .B1(n13690), .B2(n13627), .A(n582), .ZN(n6363) );
  OAI21_X2 U11370 ( .B1(n13687), .B2(n13627), .A(n583), .ZN(n6364) );
  OAI21_X2 U11371 ( .B1(n13684), .B2(n13626), .A(n584), .ZN(n6365) );
  OAI21_X2 U11372 ( .B1(n13681), .B2(n13627), .A(n585), .ZN(n6366) );
  OAI21_X2 U11373 ( .B1(n13675), .B2(n13627), .A(n587), .ZN(n6367) );
  OAI21_X2 U11374 ( .B1(n13672), .B2(n13627), .A(n588), .ZN(n6368) );
  OAI21_X2 U11375 ( .B1(n13669), .B2(n13627), .A(n589), .ZN(n6369) );
  OAI21_X2 U11376 ( .B1(n13666), .B2(n13627), .A(n590), .ZN(n6370) );
  OAI21_X2 U11377 ( .B1(n13663), .B2(n13626), .A(n591), .ZN(n6371) );
  OAI21_X2 U11378 ( .B1(n13660), .B2(n13626), .A(n592), .ZN(n6372) );
  OAI21_X2 U11379 ( .B1(n13657), .B2(n13626), .A(n593), .ZN(n6373) );
  OAI21_X2 U11380 ( .B1(n13654), .B2(n13625), .A(n594), .ZN(n6374) );
  OAI21_X2 U11381 ( .B1(n13651), .B2(n13625), .A(n595), .ZN(n6375) );
  OAI21_X2 U11382 ( .B1(n13648), .B2(n13625), .A(n596), .ZN(n6376) );
  OAI21_X2 U11383 ( .B1(n13743), .B2(n13625), .A(n566), .ZN(n6377) );
  OAI21_X2 U11384 ( .B1(n13735), .B2(n13625), .A(n567), .ZN(n6378) );
  OAI21_X2 U11385 ( .B1(n13732), .B2(n13625), .A(n568), .ZN(n6379) );
  OAI21_X2 U11386 ( .B1(n13729), .B2(n13625), .A(n569), .ZN(n6380) );
  OAI21_X2 U11387 ( .B1(n13726), .B2(n13625), .A(n570), .ZN(n6381) );
  OAI21_X2 U11388 ( .B1(n13723), .B2(n13625), .A(n571), .ZN(n6382) );
  OAI21_X2 U11389 ( .B1(n13720), .B2(n13625), .A(n572), .ZN(n6383) );
  OAI21_X2 U11390 ( .B1(n13711), .B2(n13626), .A(n575), .ZN(n6384) );
  OAI21_X2 U11391 ( .B1(n13678), .B2(n13627), .A(n586), .ZN(n6385) );
  OAI21_X2 U11392 ( .B1(n13645), .B2(n13625), .A(n597), .ZN(n6386) );
  OAI21_X2 U11393 ( .B1(n13717), .B2(n13635), .A(n504), .ZN(n6419) );
  OAI21_X2 U11394 ( .B1(n13714), .B2(n13636), .A(n505), .ZN(n6420) );
  OAI21_X2 U11395 ( .B1(n13708), .B2(n13636), .A(n507), .ZN(n6421) );
  OAI21_X2 U11396 ( .B1(n13705), .B2(n13636), .A(n508), .ZN(n6422) );
  OAI21_X2 U11397 ( .B1(n13702), .B2(n13636), .A(n509), .ZN(n6423) );
  OAI21_X2 U11398 ( .B1(n13699), .B2(n13636), .A(n510), .ZN(n6424) );
  OAI21_X2 U11399 ( .B1(n13696), .B2(n13636), .A(n511), .ZN(n6425) );
  OAI21_X2 U11400 ( .B1(n13693), .B2(n13636), .A(n512), .ZN(n6426) );
  OAI21_X2 U11401 ( .B1(n13690), .B2(n13637), .A(n513), .ZN(n6427) );
  OAI21_X2 U11402 ( .B1(n13687), .B2(n13637), .A(n514), .ZN(n6428) );
  OAI21_X2 U11403 ( .B1(n13684), .B2(n13636), .A(n515), .ZN(n6429) );
  OAI21_X2 U11404 ( .B1(n13681), .B2(n13637), .A(n516), .ZN(n6430) );
  OAI21_X2 U11405 ( .B1(n13675), .B2(n13637), .A(n518), .ZN(n6431) );
  OAI21_X2 U11406 ( .B1(n13672), .B2(n13637), .A(n519), .ZN(n6432) );
  OAI21_X2 U11407 ( .B1(n13669), .B2(n13637), .A(n520), .ZN(n6433) );
  OAI21_X2 U11408 ( .B1(n13666), .B2(n13637), .A(n521), .ZN(n6434) );
  OAI21_X2 U11409 ( .B1(n13663), .B2(n13636), .A(n522), .ZN(n6435) );
  OAI21_X2 U11410 ( .B1(n13660), .B2(n13636), .A(n523), .ZN(n6436) );
  OAI21_X2 U11411 ( .B1(n13657), .B2(n13636), .A(n524), .ZN(n6437) );
  OAI21_X2 U11412 ( .B1(n13654), .B2(n13635), .A(n525), .ZN(n6438) );
  OAI21_X2 U11413 ( .B1(n13651), .B2(n13635), .A(n526), .ZN(n6439) );
  OAI21_X2 U11414 ( .B1(n13648), .B2(n13635), .A(n527), .ZN(n6440) );
  OAI21_X2 U11415 ( .B1(n13743), .B2(n13635), .A(n497), .ZN(n6441) );
  OAI21_X2 U11416 ( .B1(n13735), .B2(n13635), .A(n498), .ZN(n6442) );
  OAI21_X2 U11417 ( .B1(n13732), .B2(n13635), .A(n499), .ZN(n6443) );
  OAI21_X2 U11418 ( .B1(n13729), .B2(n13635), .A(n500), .ZN(n6444) );
  OAI21_X2 U11419 ( .B1(n13726), .B2(n13635), .A(n501), .ZN(n6445) );
  OAI21_X2 U11420 ( .B1(n13723), .B2(n13635), .A(n502), .ZN(n6446) );
  OAI21_X2 U11421 ( .B1(n13720), .B2(n13635), .A(n503), .ZN(n6447) );
  OAI21_X2 U11422 ( .B1(n13711), .B2(n13636), .A(n506), .ZN(n6448) );
  OAI21_X2 U11423 ( .B1(n13678), .B2(n13637), .A(n517), .ZN(n6449) );
  OAI21_X2 U11424 ( .B1(n13645), .B2(n13635), .A(n528), .ZN(n6450) );
  OAI21_X2 U11425 ( .B1(n13717), .B2(n13738), .A(n411), .ZN(n6483) );
  OAI21_X2 U11426 ( .B1(n13714), .B2(n13739), .A(n413), .ZN(n6484) );
  OAI21_X2 U11427 ( .B1(n13708), .B2(n13739), .A(n417), .ZN(n6485) );
  OAI21_X2 U11428 ( .B1(n13705), .B2(n13739), .A(n419), .ZN(n6486) );
  OAI21_X2 U11429 ( .B1(n13702), .B2(n13739), .A(n421), .ZN(n6487) );
  OAI21_X2 U11430 ( .B1(n13699), .B2(n13739), .A(n423), .ZN(n6488) );
  OAI21_X2 U11431 ( .B1(n13696), .B2(n13739), .A(n425), .ZN(n6489) );
  OAI21_X2 U11432 ( .B1(n13693), .B2(n13739), .A(n427), .ZN(n6490) );
  OAI21_X2 U11433 ( .B1(n13690), .B2(n13740), .A(n429), .ZN(n6491) );
  OAI21_X2 U11434 ( .B1(n13687), .B2(n13740), .A(n431), .ZN(n6492) );
  OAI21_X2 U11435 ( .B1(n13684), .B2(n13739), .A(n433), .ZN(n6493) );
  OAI21_X2 U11436 ( .B1(n13681), .B2(n13740), .A(n435), .ZN(n6494) );
  OAI21_X2 U11437 ( .B1(n13675), .B2(n13740), .A(n439), .ZN(n6495) );
  OAI21_X2 U11438 ( .B1(n13672), .B2(n13740), .A(n441), .ZN(n6496) );
  OAI21_X2 U11439 ( .B1(n13669), .B2(n13740), .A(n443), .ZN(n6497) );
  OAI21_X2 U11440 ( .B1(n13666), .B2(n13740), .A(n445), .ZN(n6498) );
  OAI21_X2 U11441 ( .B1(n13663), .B2(n13739), .A(n447), .ZN(n6499) );
  OAI21_X2 U11442 ( .B1(n13660), .B2(n13739), .A(n449), .ZN(n6500) );
  OAI21_X2 U11443 ( .B1(n13657), .B2(n13739), .A(n451), .ZN(n6501) );
  OAI21_X2 U11444 ( .B1(n13654), .B2(n13738), .A(n453), .ZN(n6502) );
  OAI21_X2 U11445 ( .B1(n13651), .B2(n13738), .A(n455), .ZN(n6503) );
  OAI21_X2 U11446 ( .B1(n13648), .B2(n13738), .A(n457), .ZN(n6504) );
  OAI21_X2 U11447 ( .B1(n13743), .B2(n13738), .A(n397), .ZN(n6505) );
  OAI21_X2 U11448 ( .B1(n13735), .B2(n13738), .A(n399), .ZN(n6506) );
  OAI21_X2 U11449 ( .B1(n13732), .B2(n13738), .A(n401), .ZN(n6507) );
  OAI21_X2 U11450 ( .B1(n13729), .B2(n13738), .A(n403), .ZN(n6508) );
  OAI21_X2 U11451 ( .B1(n13726), .B2(n13738), .A(n405), .ZN(n6509) );
  OAI21_X2 U11452 ( .B1(n13723), .B2(n13738), .A(n407), .ZN(n6510) );
  OAI21_X2 U11453 ( .B1(n13720), .B2(n13738), .A(n409), .ZN(n6511) );
  OAI21_X2 U11454 ( .B1(n13711), .B2(n13739), .A(n415), .ZN(n6512) );
  OAI21_X2 U11455 ( .B1(n13678), .B2(n13740), .A(n437), .ZN(n6513) );
  OAI21_X2 U11456 ( .B1(n13645), .B2(n13738), .A(n459), .ZN(n6514) );
  OAI21_X2 U11457 ( .B1(n410), .B2(n13500), .A(n1412), .ZN(n6547) );
  OAI21_X2 U11458 ( .B1(n412), .B2(n13501), .A(n1413), .ZN(n6548) );
  OAI21_X2 U11459 ( .B1(n416), .B2(n13501), .A(n1415), .ZN(n6549) );
  OAI21_X2 U11460 ( .B1(n418), .B2(n13501), .A(n1416), .ZN(n6550) );
  OAI21_X2 U11461 ( .B1(n420), .B2(n13501), .A(n1417), .ZN(n6551) );
  OAI21_X2 U11462 ( .B1(n422), .B2(n13501), .A(n1418), .ZN(n6552) );
  OAI21_X2 U11463 ( .B1(n424), .B2(n13501), .A(n1419), .ZN(n6553) );
  OAI21_X2 U11464 ( .B1(n426), .B2(n13501), .A(n1420), .ZN(n6554) );
  OAI21_X2 U11465 ( .B1(n428), .B2(n13502), .A(n1421), .ZN(n6555) );
  OAI21_X2 U11466 ( .B1(n430), .B2(n13502), .A(n1422), .ZN(n6556) );
  OAI21_X2 U11467 ( .B1(n432), .B2(n13501), .A(n1423), .ZN(n6557) );
  OAI21_X2 U11468 ( .B1(n434), .B2(n13502), .A(n1424), .ZN(n6558) );
  OAI21_X2 U11469 ( .B1(n438), .B2(n13502), .A(n1426), .ZN(n6559) );
  OAI21_X2 U11470 ( .B1(n440), .B2(n13502), .A(n1427), .ZN(n6560) );
  OAI21_X2 U11471 ( .B1(n442), .B2(n13502), .A(n1428), .ZN(n6561) );
  OAI21_X2 U11472 ( .B1(n444), .B2(n13502), .A(n1429), .ZN(n6562) );
  OAI21_X2 U11473 ( .B1(n446), .B2(n13501), .A(n1430), .ZN(n6563) );
  OAI21_X2 U11474 ( .B1(n448), .B2(n13501), .A(n1431), .ZN(n6564) );
  OAI21_X2 U11475 ( .B1(n450), .B2(n13501), .A(n1432), .ZN(n6565) );
  OAI21_X2 U11476 ( .B1(n452), .B2(n13500), .A(n1433), .ZN(n6566) );
  OAI21_X2 U11477 ( .B1(n454), .B2(n13500), .A(n1434), .ZN(n6567) );
  OAI21_X2 U11478 ( .B1(n456), .B2(n13500), .A(n1435), .ZN(n6568) );
  OAI21_X2 U11479 ( .B1(n395), .B2(n13500), .A(n1405), .ZN(n6569) );
  OAI21_X2 U11480 ( .B1(n398), .B2(n13500), .A(n1406), .ZN(n6570) );
  OAI21_X2 U11481 ( .B1(n400), .B2(n13500), .A(n1407), .ZN(n6571) );
  OAI21_X2 U11482 ( .B1(n402), .B2(n13500), .A(n1408), .ZN(n6572) );
  OAI21_X2 U11483 ( .B1(n404), .B2(n13500), .A(n1409), .ZN(n6573) );
  OAI21_X2 U11484 ( .B1(n406), .B2(n13500), .A(n1410), .ZN(n6574) );
  OAI21_X2 U11485 ( .B1(n408), .B2(n13500), .A(n1411), .ZN(n6575) );
  OAI21_X2 U11486 ( .B1(n414), .B2(n13501), .A(n1414), .ZN(n6576) );
  OAI21_X2 U11487 ( .B1(n436), .B2(n13502), .A(n1425), .ZN(n6577) );
  OAI21_X2 U11488 ( .B1(n458), .B2(n13500), .A(n1436), .ZN(n6578) );
  OAI21_X2 U11489 ( .B1(n410), .B2(n13510), .A(n1345), .ZN(n6611) );
  OAI21_X2 U11490 ( .B1(n412), .B2(n13511), .A(n1346), .ZN(n6612) );
  OAI21_X2 U11491 ( .B1(n416), .B2(n13511), .A(n1348), .ZN(n6613) );
  OAI21_X2 U11492 ( .B1(n418), .B2(n13511), .A(n1349), .ZN(n6614) );
  OAI21_X2 U11493 ( .B1(n420), .B2(n13511), .A(n1350), .ZN(n6615) );
  OAI21_X2 U11494 ( .B1(n422), .B2(n13511), .A(n1351), .ZN(n6616) );
  OAI21_X2 U11495 ( .B1(n424), .B2(n13511), .A(n1352), .ZN(n6617) );
  OAI21_X2 U11496 ( .B1(n426), .B2(n13511), .A(n1353), .ZN(n6618) );
  OAI21_X2 U11497 ( .B1(n428), .B2(n13512), .A(n1354), .ZN(n6619) );
  OAI21_X2 U11498 ( .B1(n430), .B2(n13512), .A(n1355), .ZN(n6620) );
  OAI21_X2 U11499 ( .B1(n432), .B2(n13511), .A(n1356), .ZN(n6621) );
  OAI21_X2 U11500 ( .B1(n434), .B2(n13512), .A(n1357), .ZN(n6622) );
  OAI21_X2 U11501 ( .B1(n438), .B2(n13512), .A(n1359), .ZN(n6623) );
  OAI21_X2 U11502 ( .B1(n440), .B2(n13512), .A(n1360), .ZN(n6624) );
  OAI21_X2 U11503 ( .B1(n442), .B2(n13512), .A(n1361), .ZN(n6625) );
  OAI21_X2 U11504 ( .B1(n444), .B2(n13512), .A(n1362), .ZN(n6626) );
  OAI21_X2 U11505 ( .B1(n446), .B2(n13511), .A(n1363), .ZN(n6627) );
  OAI21_X2 U11506 ( .B1(n448), .B2(n13511), .A(n1364), .ZN(n6628) );
  OAI21_X2 U11507 ( .B1(n450), .B2(n13511), .A(n1365), .ZN(n6629) );
  OAI21_X2 U11508 ( .B1(n452), .B2(n13510), .A(n1366), .ZN(n6630) );
  OAI21_X2 U11509 ( .B1(n454), .B2(n13510), .A(n1367), .ZN(n6631) );
  OAI21_X2 U11510 ( .B1(n456), .B2(n13510), .A(n1368), .ZN(n6632) );
  OAI21_X2 U11511 ( .B1(n395), .B2(n13510), .A(n1338), .ZN(n6633) );
  OAI21_X2 U11512 ( .B1(n398), .B2(n13510), .A(n1339), .ZN(n6634) );
  OAI21_X2 U11513 ( .B1(n400), .B2(n13510), .A(n1340), .ZN(n6635) );
  OAI21_X2 U11514 ( .B1(n402), .B2(n13510), .A(n1341), .ZN(n6636) );
  OAI21_X2 U11515 ( .B1(n404), .B2(n13510), .A(n1342), .ZN(n6637) );
  OAI21_X2 U11516 ( .B1(n406), .B2(n13510), .A(n1343), .ZN(n6638) );
  OAI21_X2 U11517 ( .B1(n408), .B2(n13510), .A(n1344), .ZN(n6639) );
  OAI21_X2 U11518 ( .B1(n414), .B2(n13511), .A(n1347), .ZN(n6640) );
  OAI21_X2 U11519 ( .B1(n436), .B2(n13512), .A(n1358), .ZN(n6641) );
  OAI21_X2 U11520 ( .B1(n458), .B2(n13510), .A(n1369), .ZN(n6642) );
  OAI21_X2 U11521 ( .B1(n410), .B2(n13520), .A(n1279), .ZN(n6675) );
  OAI21_X2 U11522 ( .B1(n412), .B2(n13521), .A(n1280), .ZN(n6676) );
  OAI21_X2 U11523 ( .B1(n416), .B2(n13521), .A(n1282), .ZN(n6677) );
  OAI21_X2 U11524 ( .B1(n418), .B2(n13521), .A(n1283), .ZN(n6678) );
  OAI21_X2 U11525 ( .B1(n420), .B2(n13521), .A(n1284), .ZN(n6679) );
  OAI21_X2 U11526 ( .B1(n422), .B2(n13521), .A(n1285), .ZN(n6680) );
  OAI21_X2 U11527 ( .B1(n424), .B2(n13521), .A(n1286), .ZN(n6681) );
  OAI21_X2 U11528 ( .B1(n426), .B2(n13521), .A(n1287), .ZN(n6682) );
  OAI21_X2 U11529 ( .B1(n428), .B2(n13522), .A(n1288), .ZN(n6683) );
  OAI21_X2 U11530 ( .B1(n430), .B2(n13522), .A(n1289), .ZN(n6684) );
  OAI21_X2 U11531 ( .B1(n432), .B2(n13521), .A(n1290), .ZN(n6685) );
  OAI21_X2 U11532 ( .B1(n434), .B2(n13522), .A(n1291), .ZN(n6686) );
  OAI21_X2 U11533 ( .B1(n438), .B2(n13522), .A(n1293), .ZN(n6687) );
  OAI21_X2 U11534 ( .B1(n440), .B2(n13522), .A(n1294), .ZN(n6688) );
  OAI21_X2 U11535 ( .B1(n442), .B2(n13522), .A(n1295), .ZN(n6689) );
  OAI21_X2 U11536 ( .B1(n444), .B2(n13522), .A(n1296), .ZN(n6690) );
  OAI21_X2 U11537 ( .B1(n446), .B2(n13521), .A(n1297), .ZN(n6691) );
  OAI21_X2 U11538 ( .B1(n448), .B2(n13521), .A(n1298), .ZN(n6692) );
  OAI21_X2 U11539 ( .B1(n450), .B2(n13521), .A(n1299), .ZN(n6693) );
  OAI21_X2 U11540 ( .B1(n452), .B2(n13520), .A(n1300), .ZN(n6694) );
  OAI21_X2 U11541 ( .B1(n454), .B2(n13520), .A(n1301), .ZN(n6695) );
  OAI21_X2 U11542 ( .B1(n456), .B2(n13520), .A(n1302), .ZN(n6696) );
  OAI21_X2 U11543 ( .B1(n395), .B2(n13520), .A(n1272), .ZN(n6697) );
  OAI21_X2 U11544 ( .B1(n398), .B2(n13520), .A(n1273), .ZN(n6698) );
  OAI21_X2 U11545 ( .B1(n400), .B2(n13520), .A(n1274), .ZN(n6699) );
  OAI21_X2 U11546 ( .B1(n402), .B2(n13520), .A(n1275), .ZN(n6700) );
  OAI21_X2 U11547 ( .B1(n404), .B2(n13520), .A(n1276), .ZN(n6701) );
  OAI21_X2 U11548 ( .B1(n406), .B2(n13520), .A(n1277), .ZN(n6702) );
  OAI21_X2 U11549 ( .B1(n408), .B2(n13520), .A(n1278), .ZN(n6703) );
  OAI21_X2 U11550 ( .B1(n414), .B2(n13521), .A(n1281), .ZN(n6704) );
  OAI21_X2 U11551 ( .B1(n436), .B2(n13522), .A(n1292), .ZN(n6705) );
  OAI21_X2 U11552 ( .B1(n458), .B2(n13520), .A(n1303), .ZN(n6706) );
  OAI21_X2 U11553 ( .B1(n13718), .B2(n13530), .A(n1211), .ZN(n6739) );
  OAI21_X2 U11554 ( .B1(n13715), .B2(n13531), .A(n1212), .ZN(n6740) );
  OAI21_X2 U11555 ( .B1(n13709), .B2(n13531), .A(n1214), .ZN(n6741) );
  OAI21_X2 U11556 ( .B1(n13706), .B2(n13531), .A(n1215), .ZN(n6742) );
  OAI21_X2 U11557 ( .B1(n13703), .B2(n13531), .A(n1216), .ZN(n6743) );
  OAI21_X2 U11558 ( .B1(n13700), .B2(n13531), .A(n1217), .ZN(n6744) );
  OAI21_X2 U11559 ( .B1(n13697), .B2(n13531), .A(n1218), .ZN(n6745) );
  OAI21_X2 U11560 ( .B1(n13694), .B2(n13531), .A(n1219), .ZN(n6746) );
  OAI21_X2 U11561 ( .B1(n13691), .B2(n13532), .A(n1220), .ZN(n6747) );
  OAI21_X2 U11562 ( .B1(n13688), .B2(n13532), .A(n1221), .ZN(n6748) );
  OAI21_X2 U11563 ( .B1(n13685), .B2(n13531), .A(n1222), .ZN(n6749) );
  OAI21_X2 U11564 ( .B1(n13682), .B2(n13532), .A(n1223), .ZN(n6750) );
  OAI21_X2 U11565 ( .B1(n13676), .B2(n13532), .A(n1225), .ZN(n6751) );
  OAI21_X2 U11566 ( .B1(n13673), .B2(n13532), .A(n1226), .ZN(n6752) );
  OAI21_X2 U11567 ( .B1(n13670), .B2(n13532), .A(n1227), .ZN(n6753) );
  OAI21_X2 U11568 ( .B1(n13667), .B2(n13532), .A(n1228), .ZN(n6754) );
  OAI21_X2 U11569 ( .B1(n13664), .B2(n13531), .A(n1229), .ZN(n6755) );
  OAI21_X2 U11570 ( .B1(n13661), .B2(n13531), .A(n1230), .ZN(n6756) );
  OAI21_X2 U11571 ( .B1(n13658), .B2(n13531), .A(n1231), .ZN(n6757) );
  OAI21_X2 U11572 ( .B1(n13655), .B2(n13530), .A(n1232), .ZN(n6758) );
  OAI21_X2 U11573 ( .B1(n13652), .B2(n13530), .A(n1233), .ZN(n6759) );
  OAI21_X2 U11574 ( .B1(n13649), .B2(n13530), .A(n1234), .ZN(n6760) );
  OAI21_X2 U11575 ( .B1(n13744), .B2(n13530), .A(n1204), .ZN(n6761) );
  OAI21_X2 U11576 ( .B1(n13736), .B2(n13530), .A(n1205), .ZN(n6762) );
  OAI21_X2 U11577 ( .B1(n13733), .B2(n13530), .A(n1206), .ZN(n6763) );
  OAI21_X2 U11578 ( .B1(n13730), .B2(n13530), .A(n1207), .ZN(n6764) );
  OAI21_X2 U11579 ( .B1(n13727), .B2(n13530), .A(n1208), .ZN(n6765) );
  OAI21_X2 U11580 ( .B1(n13724), .B2(n13530), .A(n1209), .ZN(n6766) );
  OAI21_X2 U11581 ( .B1(n13721), .B2(n13530), .A(n1210), .ZN(n6767) );
  OAI21_X2 U11582 ( .B1(n13712), .B2(n13531), .A(n1213), .ZN(n6768) );
  OAI21_X2 U11583 ( .B1(n13679), .B2(n13532), .A(n1224), .ZN(n6769) );
  OAI21_X2 U11584 ( .B1(n13646), .B2(n13530), .A(n1235), .ZN(n6770) );
  OAI21_X2 U11585 ( .B1(n13718), .B2(n13540), .A(n1144), .ZN(n6803) );
  OAI21_X2 U11586 ( .B1(n13715), .B2(n13541), .A(n1145), .ZN(n6804) );
  OAI21_X2 U11587 ( .B1(n13709), .B2(n13541), .A(n1147), .ZN(n6805) );
  OAI21_X2 U11588 ( .B1(n13706), .B2(n13541), .A(n1148), .ZN(n6806) );
  OAI21_X2 U11589 ( .B1(n13703), .B2(n13541), .A(n1149), .ZN(n6807) );
  OAI21_X2 U11590 ( .B1(n13700), .B2(n13541), .A(n1150), .ZN(n6808) );
  OAI21_X2 U11591 ( .B1(n13697), .B2(n13541), .A(n1151), .ZN(n6809) );
  OAI21_X2 U11592 ( .B1(n13694), .B2(n13541), .A(n1152), .ZN(n6810) );
  OAI21_X2 U11593 ( .B1(n13691), .B2(n13542), .A(n1153), .ZN(n6811) );
  OAI21_X2 U11594 ( .B1(n13688), .B2(n13542), .A(n1154), .ZN(n6812) );
  OAI21_X2 U11595 ( .B1(n13685), .B2(n13541), .A(n1155), .ZN(n6813) );
  OAI21_X2 U11596 ( .B1(n13682), .B2(n13542), .A(n1156), .ZN(n6814) );
  OAI21_X2 U11597 ( .B1(n13676), .B2(n13542), .A(n1158), .ZN(n6815) );
  OAI21_X2 U11598 ( .B1(n13673), .B2(n13542), .A(n1159), .ZN(n6816) );
  OAI21_X2 U11599 ( .B1(n13670), .B2(n13542), .A(n1160), .ZN(n6817) );
  OAI21_X2 U11600 ( .B1(n13667), .B2(n13542), .A(n1161), .ZN(n6818) );
  OAI21_X2 U11601 ( .B1(n13664), .B2(n13541), .A(n1162), .ZN(n6819) );
  OAI21_X2 U11602 ( .B1(n13661), .B2(n13541), .A(n1163), .ZN(n6820) );
  OAI21_X2 U11603 ( .B1(n13658), .B2(n13541), .A(n1164), .ZN(n6821) );
  OAI21_X2 U11604 ( .B1(n13655), .B2(n13540), .A(n1165), .ZN(n6822) );
  OAI21_X2 U11605 ( .B1(n13652), .B2(n13540), .A(n1166), .ZN(n6823) );
  OAI21_X2 U11606 ( .B1(n13649), .B2(n13540), .A(n1167), .ZN(n6824) );
  OAI21_X2 U11607 ( .B1(n13744), .B2(n13540), .A(n1137), .ZN(n6825) );
  OAI21_X2 U11608 ( .B1(n13736), .B2(n13540), .A(n1138), .ZN(n6826) );
  OAI21_X2 U11609 ( .B1(n13733), .B2(n13540), .A(n1139), .ZN(n6827) );
  OAI21_X2 U11610 ( .B1(n13730), .B2(n13540), .A(n1140), .ZN(n6828) );
  OAI21_X2 U11611 ( .B1(n13727), .B2(n13540), .A(n1141), .ZN(n6829) );
  OAI21_X2 U11612 ( .B1(n13724), .B2(n13540), .A(n1142), .ZN(n6830) );
  OAI21_X2 U11613 ( .B1(n13721), .B2(n13540), .A(n1143), .ZN(n6831) );
  OAI21_X2 U11614 ( .B1(n13712), .B2(n13541), .A(n1146), .ZN(n6832) );
  OAI21_X2 U11615 ( .B1(n13679), .B2(n13542), .A(n1157), .ZN(n6833) );
  OAI21_X2 U11616 ( .B1(n13646), .B2(n13540), .A(n1168), .ZN(n6834) );
  OAI21_X2 U11617 ( .B1(n13718), .B2(n13555), .A(n1045), .ZN(n6867) );
  OAI21_X2 U11618 ( .B1(n13715), .B2(n13556), .A(n1046), .ZN(n6868) );
  OAI21_X2 U11619 ( .B1(n13709), .B2(n13556), .A(n1048), .ZN(n6869) );
  OAI21_X2 U11620 ( .B1(n13706), .B2(n13556), .A(n1049), .ZN(n6870) );
  OAI21_X2 U11621 ( .B1(n13703), .B2(n13556), .A(n1050), .ZN(n6871) );
  OAI21_X2 U11622 ( .B1(n13700), .B2(n13556), .A(n1051), .ZN(n6872) );
  OAI21_X2 U11623 ( .B1(n13697), .B2(n13556), .A(n1052), .ZN(n6873) );
  OAI21_X2 U11624 ( .B1(n13694), .B2(n13556), .A(n1053), .ZN(n6874) );
  OAI21_X2 U11625 ( .B1(n13691), .B2(n13557), .A(n1054), .ZN(n6875) );
  OAI21_X2 U11626 ( .B1(n13688), .B2(n13557), .A(n1055), .ZN(n6876) );
  OAI21_X2 U11627 ( .B1(n13685), .B2(n13556), .A(n1056), .ZN(n6877) );
  OAI21_X2 U11628 ( .B1(n13682), .B2(n13557), .A(n1057), .ZN(n6878) );
  OAI21_X2 U11629 ( .B1(n13676), .B2(n13557), .A(n1059), .ZN(n6879) );
  OAI21_X2 U11630 ( .B1(n13673), .B2(n13557), .A(n1060), .ZN(n6880) );
  OAI21_X2 U11631 ( .B1(n13670), .B2(n13557), .A(n1061), .ZN(n6881) );
  OAI21_X2 U11632 ( .B1(n13667), .B2(n13557), .A(n1062), .ZN(n6882) );
  OAI21_X2 U11633 ( .B1(n13664), .B2(n13556), .A(n1063), .ZN(n6883) );
  OAI21_X2 U11634 ( .B1(n13661), .B2(n13556), .A(n1064), .ZN(n6884) );
  OAI21_X2 U11635 ( .B1(n13658), .B2(n13556), .A(n1065), .ZN(n6885) );
  OAI21_X2 U11636 ( .B1(n13655), .B2(n13555), .A(n1066), .ZN(n6886) );
  OAI21_X2 U11637 ( .B1(n13652), .B2(n13555), .A(n1067), .ZN(n6887) );
  OAI21_X2 U11638 ( .B1(n13649), .B2(n13555), .A(n1068), .ZN(n6888) );
  OAI21_X2 U11639 ( .B1(n13744), .B2(n13555), .A(n1038), .ZN(n6889) );
  OAI21_X2 U11640 ( .B1(n13736), .B2(n13555), .A(n1039), .ZN(n6890) );
  OAI21_X2 U11641 ( .B1(n13733), .B2(n13555), .A(n1040), .ZN(n6891) );
  OAI21_X2 U11642 ( .B1(n13730), .B2(n13555), .A(n1041), .ZN(n6892) );
  OAI21_X2 U11643 ( .B1(n13727), .B2(n13555), .A(n1042), .ZN(n6893) );
  OAI21_X2 U11644 ( .B1(n13724), .B2(n13555), .A(n1043), .ZN(n6894) );
  OAI21_X2 U11645 ( .B1(n13721), .B2(n13555), .A(n1044), .ZN(n6895) );
  OAI21_X2 U11646 ( .B1(n13712), .B2(n13556), .A(n1047), .ZN(n6896) );
  OAI21_X2 U11647 ( .B1(n13679), .B2(n13557), .A(n1058), .ZN(n6897) );
  OAI21_X2 U11648 ( .B1(n13646), .B2(n13555), .A(n1069), .ZN(n6898) );
  OAI21_X2 U11649 ( .B1(n13718), .B2(n13565), .A(n978), .ZN(n6931) );
  OAI21_X2 U11650 ( .B1(n13715), .B2(n13566), .A(n979), .ZN(n6932) );
  OAI21_X2 U11651 ( .B1(n13709), .B2(n13566), .A(n981), .ZN(n6933) );
  OAI21_X2 U11652 ( .B1(n13706), .B2(n13566), .A(n982), .ZN(n6934) );
  OAI21_X2 U11653 ( .B1(n13703), .B2(n13566), .A(n983), .ZN(n6935) );
  OAI21_X2 U11654 ( .B1(n13700), .B2(n13566), .A(n984), .ZN(n6936) );
  OAI21_X2 U11655 ( .B1(n13697), .B2(n13566), .A(n985), .ZN(n6937) );
  OAI21_X2 U11656 ( .B1(n13694), .B2(n13566), .A(n986), .ZN(n6938) );
  OAI21_X2 U11657 ( .B1(n13691), .B2(n13567), .A(n987), .ZN(n6939) );
  OAI21_X2 U11658 ( .B1(n13688), .B2(n13567), .A(n988), .ZN(n6940) );
  OAI21_X2 U11659 ( .B1(n13685), .B2(n13566), .A(n989), .ZN(n6941) );
  OAI21_X2 U11660 ( .B1(n13682), .B2(n13567), .A(n990), .ZN(n6942) );
  OAI21_X2 U11661 ( .B1(n13676), .B2(n13567), .A(n992), .ZN(n6943) );
  OAI21_X2 U11662 ( .B1(n13673), .B2(n13567), .A(n993), .ZN(n6944) );
  OAI21_X2 U11663 ( .B1(n13670), .B2(n13567), .A(n994), .ZN(n6945) );
  OAI21_X2 U11664 ( .B1(n13667), .B2(n13567), .A(n995), .ZN(n6946) );
  OAI21_X2 U11665 ( .B1(n13664), .B2(n13566), .A(n996), .ZN(n6947) );
  OAI21_X2 U11666 ( .B1(n13661), .B2(n13566), .A(n997), .ZN(n6948) );
  OAI21_X2 U11667 ( .B1(n13658), .B2(n13566), .A(n998), .ZN(n6949) );
  OAI21_X2 U11668 ( .B1(n13655), .B2(n13565), .A(n999), .ZN(n6950) );
  OAI21_X2 U11669 ( .B1(n13652), .B2(n13565), .A(n1000), .ZN(n6951) );
  OAI21_X2 U11670 ( .B1(n13649), .B2(n13565), .A(n1001), .ZN(n6952) );
  OAI21_X2 U11671 ( .B1(n13744), .B2(n13565), .A(n971), .ZN(n6953) );
  OAI21_X2 U11672 ( .B1(n13736), .B2(n13565), .A(n972), .ZN(n6954) );
  OAI21_X2 U11673 ( .B1(n13733), .B2(n13565), .A(n973), .ZN(n6955) );
  OAI21_X2 U11674 ( .B1(n13730), .B2(n13565), .A(n974), .ZN(n6956) );
  OAI21_X2 U11675 ( .B1(n13727), .B2(n13565), .A(n975), .ZN(n6957) );
  OAI21_X2 U11676 ( .B1(n13724), .B2(n13565), .A(n976), .ZN(n6958) );
  OAI21_X2 U11677 ( .B1(n13721), .B2(n13565), .A(n977), .ZN(n6959) );
  OAI21_X2 U11678 ( .B1(n13712), .B2(n13566), .A(n980), .ZN(n6960) );
  OAI21_X2 U11679 ( .B1(n13679), .B2(n13567), .A(n991), .ZN(n6961) );
  OAI21_X2 U11680 ( .B1(n13646), .B2(n13565), .A(n1002), .ZN(n6962) );
  OAI21_X2 U11681 ( .B1(n13718), .B2(n13575), .A(n912), .ZN(n6995) );
  OAI21_X2 U11682 ( .B1(n13715), .B2(n13576), .A(n913), .ZN(n6996) );
  OAI21_X2 U11683 ( .B1(n13709), .B2(n13576), .A(n915), .ZN(n6997) );
  OAI21_X2 U11684 ( .B1(n13706), .B2(n13576), .A(n916), .ZN(n6998) );
  OAI21_X2 U11685 ( .B1(n13703), .B2(n13576), .A(n917), .ZN(n6999) );
  OAI21_X2 U11686 ( .B1(n13700), .B2(n13576), .A(n918), .ZN(n7000) );
  OAI21_X2 U11687 ( .B1(n13697), .B2(n13576), .A(n919), .ZN(n7001) );
  OAI21_X2 U11688 ( .B1(n13694), .B2(n13576), .A(n920), .ZN(n7002) );
  OAI21_X2 U11689 ( .B1(n13691), .B2(n13577), .A(n921), .ZN(n7003) );
  OAI21_X2 U11690 ( .B1(n13688), .B2(n13577), .A(n922), .ZN(n7004) );
  OAI21_X2 U11691 ( .B1(n13685), .B2(n13576), .A(n923), .ZN(n7005) );
  OAI21_X2 U11692 ( .B1(n13682), .B2(n13577), .A(n924), .ZN(n7006) );
  OAI21_X2 U11693 ( .B1(n13676), .B2(n13577), .A(n926), .ZN(n7007) );
  OAI21_X2 U11694 ( .B1(n13673), .B2(n13577), .A(n927), .ZN(n7008) );
  OAI21_X2 U11695 ( .B1(n13670), .B2(n13577), .A(n928), .ZN(n7009) );
  OAI21_X2 U11696 ( .B1(n13667), .B2(n13577), .A(n929), .ZN(n7010) );
  OAI21_X2 U11697 ( .B1(n13664), .B2(n13576), .A(n930), .ZN(n7011) );
  OAI21_X2 U11698 ( .B1(n13661), .B2(n13576), .A(n931), .ZN(n7012) );
  OAI21_X2 U11699 ( .B1(n13658), .B2(n13576), .A(n932), .ZN(n7013) );
  OAI21_X2 U11700 ( .B1(n13655), .B2(n13575), .A(n933), .ZN(n7014) );
  OAI21_X2 U11701 ( .B1(n13652), .B2(n13575), .A(n934), .ZN(n7015) );
  OAI21_X2 U11702 ( .B1(n13649), .B2(n13575), .A(n935), .ZN(n7016) );
  OAI21_X2 U11703 ( .B1(n13744), .B2(n13575), .A(n905), .ZN(n7017) );
  OAI21_X2 U11704 ( .B1(n13736), .B2(n13575), .A(n906), .ZN(n7018) );
  OAI21_X2 U11705 ( .B1(n13733), .B2(n13575), .A(n907), .ZN(n7019) );
  OAI21_X2 U11706 ( .B1(n13730), .B2(n13575), .A(n908), .ZN(n7020) );
  OAI21_X2 U11707 ( .B1(n13727), .B2(n13575), .A(n909), .ZN(n7021) );
  OAI21_X2 U11708 ( .B1(n13724), .B2(n13575), .A(n910), .ZN(n7022) );
  OAI21_X2 U11709 ( .B1(n13721), .B2(n13575), .A(n911), .ZN(n7023) );
  OAI21_X2 U11710 ( .B1(n13712), .B2(n13576), .A(n914), .ZN(n7024) );
  OAI21_X2 U11711 ( .B1(n13679), .B2(n13577), .A(n925), .ZN(n7025) );
  OAI21_X2 U11712 ( .B1(n13646), .B2(n13575), .A(n936), .ZN(n7026) );
  OAI21_X2 U11713 ( .B1(n13718), .B2(n13585), .A(n845), .ZN(n7059) );
  OAI21_X2 U11714 ( .B1(n13715), .B2(n13586), .A(n846), .ZN(n7060) );
  OAI21_X2 U11715 ( .B1(n13709), .B2(n13586), .A(n848), .ZN(n7061) );
  OAI21_X2 U11716 ( .B1(n13706), .B2(n13586), .A(n849), .ZN(n7062) );
  OAI21_X2 U11717 ( .B1(n13703), .B2(n13586), .A(n850), .ZN(n7063) );
  OAI21_X2 U11718 ( .B1(n13700), .B2(n13586), .A(n851), .ZN(n7064) );
  OAI21_X2 U11719 ( .B1(n13697), .B2(n13586), .A(n852), .ZN(n7065) );
  OAI21_X2 U11720 ( .B1(n13694), .B2(n13586), .A(n853), .ZN(n7066) );
  OAI21_X2 U11721 ( .B1(n13691), .B2(n13587), .A(n854), .ZN(n7067) );
  OAI21_X2 U11722 ( .B1(n13688), .B2(n13587), .A(n855), .ZN(n7068) );
  OAI21_X2 U11723 ( .B1(n13685), .B2(n13586), .A(n856), .ZN(n7069) );
  OAI21_X2 U11724 ( .B1(n13682), .B2(n13587), .A(n857), .ZN(n7070) );
  OAI21_X2 U11725 ( .B1(n13676), .B2(n13587), .A(n859), .ZN(n7071) );
  OAI21_X2 U11726 ( .B1(n13673), .B2(n13587), .A(n860), .ZN(n7072) );
  OAI21_X2 U11727 ( .B1(n13670), .B2(n13587), .A(n861), .ZN(n7073) );
  OAI21_X2 U11728 ( .B1(n13667), .B2(n13587), .A(n862), .ZN(n7074) );
  OAI21_X2 U11729 ( .B1(n13664), .B2(n13586), .A(n863), .ZN(n7075) );
  OAI21_X2 U11730 ( .B1(n13661), .B2(n13586), .A(n864), .ZN(n7076) );
  OAI21_X2 U11731 ( .B1(n13658), .B2(n13586), .A(n865), .ZN(n7077) );
  OAI21_X2 U11732 ( .B1(n13655), .B2(n13585), .A(n866), .ZN(n7078) );
  OAI21_X2 U11733 ( .B1(n13652), .B2(n13585), .A(n867), .ZN(n7079) );
  OAI21_X2 U11734 ( .B1(n13649), .B2(n13585), .A(n868), .ZN(n7080) );
  OAI21_X2 U11735 ( .B1(n13744), .B2(n13585), .A(n838), .ZN(n7081) );
  OAI21_X2 U11736 ( .B1(n13736), .B2(n13585), .A(n839), .ZN(n7082) );
  OAI21_X2 U11737 ( .B1(n13733), .B2(n13585), .A(n840), .ZN(n7083) );
  OAI21_X2 U11738 ( .B1(n13730), .B2(n13585), .A(n841), .ZN(n7084) );
  OAI21_X2 U11739 ( .B1(n13727), .B2(n13585), .A(n842), .ZN(n7085) );
  OAI21_X2 U11740 ( .B1(n13724), .B2(n13585), .A(n843), .ZN(n7086) );
  OAI21_X2 U11741 ( .B1(n13721), .B2(n13585), .A(n844), .ZN(n7087) );
  OAI21_X2 U11742 ( .B1(n13712), .B2(n13586), .A(n847), .ZN(n7088) );
  OAI21_X2 U11743 ( .B1(n13679), .B2(n13587), .A(n858), .ZN(n7089) );
  OAI21_X2 U11744 ( .B1(n13646), .B2(n13585), .A(n869), .ZN(n7090) );
  OAI21_X2 U11745 ( .B1(n13717), .B2(n13595), .A(n775), .ZN(n7123) );
  OAI21_X2 U11746 ( .B1(n13714), .B2(n13596), .A(n776), .ZN(n7124) );
  OAI21_X2 U11747 ( .B1(n13708), .B2(n13596), .A(n778), .ZN(n7125) );
  OAI21_X2 U11748 ( .B1(n13705), .B2(n13596), .A(n779), .ZN(n7126) );
  OAI21_X2 U11749 ( .B1(n13702), .B2(n13596), .A(n780), .ZN(n7127) );
  OAI21_X2 U11750 ( .B1(n13699), .B2(n13596), .A(n781), .ZN(n7128) );
  OAI21_X2 U11751 ( .B1(n13696), .B2(n13596), .A(n782), .ZN(n7129) );
  OAI21_X2 U11752 ( .B1(n13693), .B2(n13596), .A(n783), .ZN(n7130) );
  OAI21_X2 U11753 ( .B1(n13690), .B2(n13597), .A(n784), .ZN(n7131) );
  OAI21_X2 U11754 ( .B1(n13687), .B2(n13597), .A(n785), .ZN(n7132) );
  OAI21_X2 U11755 ( .B1(n13684), .B2(n13596), .A(n786), .ZN(n7133) );
  OAI21_X2 U11756 ( .B1(n13681), .B2(n13597), .A(n787), .ZN(n7134) );
  OAI21_X2 U11757 ( .B1(n13675), .B2(n13597), .A(n789), .ZN(n7135) );
  OAI21_X2 U11758 ( .B1(n13672), .B2(n13597), .A(n790), .ZN(n7136) );
  OAI21_X2 U11759 ( .B1(n13669), .B2(n13597), .A(n791), .ZN(n7137) );
  OAI21_X2 U11760 ( .B1(n13666), .B2(n13597), .A(n792), .ZN(n7138) );
  OAI21_X2 U11761 ( .B1(n13663), .B2(n13596), .A(n793), .ZN(n7139) );
  OAI21_X2 U11762 ( .B1(n13660), .B2(n13596), .A(n794), .ZN(n7140) );
  OAI21_X2 U11763 ( .B1(n13657), .B2(n13596), .A(n795), .ZN(n7141) );
  OAI21_X2 U11764 ( .B1(n13654), .B2(n13595), .A(n796), .ZN(n7142) );
  OAI21_X2 U11765 ( .B1(n13651), .B2(n13595), .A(n797), .ZN(n7143) );
  OAI21_X2 U11766 ( .B1(n13648), .B2(n13595), .A(n798), .ZN(n7144) );
  OAI21_X2 U11767 ( .B1(n13743), .B2(n13595), .A(n768), .ZN(n7145) );
  OAI21_X2 U11768 ( .B1(n13735), .B2(n13595), .A(n769), .ZN(n7146) );
  OAI21_X2 U11769 ( .B1(n13732), .B2(n13595), .A(n770), .ZN(n7147) );
  OAI21_X2 U11770 ( .B1(n13729), .B2(n13595), .A(n771), .ZN(n7148) );
  OAI21_X2 U11771 ( .B1(n13726), .B2(n13595), .A(n772), .ZN(n7149) );
  OAI21_X2 U11772 ( .B1(n13723), .B2(n13595), .A(n773), .ZN(n7150) );
  OAI21_X2 U11773 ( .B1(n13720), .B2(n13595), .A(n774), .ZN(n7151) );
  OAI21_X2 U11774 ( .B1(n13711), .B2(n13596), .A(n777), .ZN(n7152) );
  OAI21_X2 U11775 ( .B1(n13678), .B2(n13597), .A(n788), .ZN(n7153) );
  OAI21_X2 U11776 ( .B1(n13645), .B2(n13595), .A(n799), .ZN(n7154) );
  OAI21_X2 U11777 ( .B1(n13717), .B2(n13610), .A(n673), .ZN(n7187) );
  OAI21_X2 U11778 ( .B1(n13714), .B2(n13611), .A(n674), .ZN(n7188) );
  OAI21_X2 U11779 ( .B1(n13708), .B2(n13611), .A(n676), .ZN(n7189) );
  OAI21_X2 U11780 ( .B1(n13705), .B2(n13611), .A(n677), .ZN(n7190) );
  OAI21_X2 U11781 ( .B1(n13702), .B2(n13611), .A(n678), .ZN(n7191) );
  OAI21_X2 U11782 ( .B1(n13699), .B2(n13611), .A(n679), .ZN(n7192) );
  OAI21_X2 U11783 ( .B1(n13696), .B2(n13611), .A(n680), .ZN(n7193) );
  OAI21_X2 U11784 ( .B1(n13693), .B2(n13611), .A(n681), .ZN(n7194) );
  OAI21_X2 U11785 ( .B1(n13690), .B2(n13612), .A(n682), .ZN(n7195) );
  OAI21_X2 U11786 ( .B1(n13687), .B2(n13612), .A(n683), .ZN(n7196) );
  OAI21_X2 U11787 ( .B1(n13684), .B2(n13611), .A(n684), .ZN(n7197) );
  OAI21_X2 U11788 ( .B1(n13681), .B2(n13612), .A(n685), .ZN(n7198) );
  OAI21_X2 U11789 ( .B1(n13675), .B2(n13612), .A(n687), .ZN(n7199) );
  OAI21_X2 U11790 ( .B1(n13672), .B2(n13612), .A(n688), .ZN(n7200) );
  OAI21_X2 U11791 ( .B1(n13669), .B2(n13612), .A(n689), .ZN(n7201) );
  OAI21_X2 U11792 ( .B1(n13666), .B2(n13612), .A(n690), .ZN(n7202) );
  OAI21_X2 U11793 ( .B1(n13663), .B2(n13611), .A(n691), .ZN(n7203) );
  OAI21_X2 U11794 ( .B1(n13660), .B2(n13611), .A(n692), .ZN(n7204) );
  OAI21_X2 U11795 ( .B1(n13657), .B2(n13611), .A(n693), .ZN(n7205) );
  OAI21_X2 U11796 ( .B1(n13654), .B2(n13610), .A(n694), .ZN(n7206) );
  OAI21_X2 U11797 ( .B1(n13651), .B2(n13610), .A(n695), .ZN(n7207) );
  OAI21_X2 U11798 ( .B1(n13648), .B2(n13610), .A(n696), .ZN(n7208) );
  OAI21_X2 U11799 ( .B1(n13743), .B2(n13610), .A(n666), .ZN(n7209) );
  OAI21_X2 U11800 ( .B1(n13735), .B2(n13610), .A(n667), .ZN(n7210) );
  OAI21_X2 U11801 ( .B1(n13732), .B2(n13610), .A(n668), .ZN(n7211) );
  OAI21_X2 U11802 ( .B1(n13729), .B2(n13610), .A(n669), .ZN(n7212) );
  OAI21_X2 U11803 ( .B1(n13726), .B2(n13610), .A(n670), .ZN(n7213) );
  OAI21_X2 U11804 ( .B1(n13723), .B2(n13610), .A(n671), .ZN(n7214) );
  OAI21_X2 U11805 ( .B1(n13720), .B2(n13610), .A(n672), .ZN(n7215) );
  OAI21_X2 U11806 ( .B1(n13711), .B2(n13611), .A(n675), .ZN(n7216) );
  OAI21_X2 U11807 ( .B1(n13678), .B2(n13612), .A(n686), .ZN(n7217) );
  OAI21_X2 U11808 ( .B1(n13645), .B2(n13610), .A(n697), .ZN(n7218) );
  OAI21_X2 U11809 ( .B1(n13458), .B2(n13285), .A(n2215), .ZN(n7251) );
  OAI21_X2 U11810 ( .B1(n13455), .B2(n13286), .A(n2216), .ZN(n7252) );
  OAI21_X2 U11811 ( .B1(n13449), .B2(n13286), .A(n2218), .ZN(n7253) );
  OAI21_X2 U11812 ( .B1(n13446), .B2(n13286), .A(n2219), .ZN(n7254) );
  OAI21_X2 U11813 ( .B1(n13443), .B2(n13286), .A(n2220), .ZN(n7255) );
  OAI21_X2 U11814 ( .B1(n13440), .B2(n13286), .A(n2221), .ZN(n7256) );
  OAI21_X2 U11815 ( .B1(n13437), .B2(n13286), .A(n2222), .ZN(n7257) );
  OAI21_X2 U11816 ( .B1(n13434), .B2(n13286), .A(n2223), .ZN(n7258) );
  OAI21_X2 U11817 ( .B1(n13431), .B2(n13287), .A(n2224), .ZN(n7259) );
  OAI21_X2 U11818 ( .B1(n13428), .B2(n13287), .A(n2225), .ZN(n7260) );
  OAI21_X2 U11819 ( .B1(n13425), .B2(n13286), .A(n2226), .ZN(n7261) );
  OAI21_X2 U11820 ( .B1(n13422), .B2(n13287), .A(n2227), .ZN(n7262) );
  OAI21_X2 U11821 ( .B1(n13416), .B2(n13287), .A(n2229), .ZN(n7263) );
  OAI21_X2 U11822 ( .B1(n13413), .B2(n13287), .A(n2230), .ZN(n7264) );
  OAI21_X2 U11823 ( .B1(n13410), .B2(n13287), .A(n2231), .ZN(n7265) );
  OAI21_X2 U11824 ( .B1(n13407), .B2(n13287), .A(n2232), .ZN(n7266) );
  OAI21_X2 U11825 ( .B1(n13404), .B2(n13286), .A(n2233), .ZN(n7267) );
  OAI21_X2 U11826 ( .B1(n13401), .B2(n13286), .A(n2234), .ZN(n7268) );
  OAI21_X2 U11827 ( .B1(n13398), .B2(n13286), .A(n2235), .ZN(n7269) );
  OAI21_X2 U11828 ( .B1(n13395), .B2(n13285), .A(n2236), .ZN(n7270) );
  OAI21_X2 U11829 ( .B1(n13392), .B2(n13285), .A(n2237), .ZN(n7271) );
  OAI21_X2 U11830 ( .B1(n13389), .B2(n13285), .A(n2238), .ZN(n7272) );
  OAI21_X2 U11831 ( .B1(n13484), .B2(n13285), .A(n2208), .ZN(n7273) );
  OAI21_X2 U11832 ( .B1(n13476), .B2(n13285), .A(n2209), .ZN(n7274) );
  OAI21_X2 U11833 ( .B1(n13473), .B2(n13285), .A(n2210), .ZN(n7275) );
  OAI21_X2 U11834 ( .B1(n13470), .B2(n13285), .A(n2211), .ZN(n7276) );
  OAI21_X2 U11835 ( .B1(n13467), .B2(n13285), .A(n2212), .ZN(n7277) );
  OAI21_X2 U11836 ( .B1(n13464), .B2(n13285), .A(n2213), .ZN(n7278) );
  OAI21_X2 U11837 ( .B1(n13461), .B2(n13285), .A(n2214), .ZN(n7279) );
  OAI21_X2 U11838 ( .B1(n13452), .B2(n13286), .A(n2217), .ZN(n7280) );
  OAI21_X2 U11839 ( .B1(n13419), .B2(n13287), .A(n2228), .ZN(n7281) );
  OAI21_X2 U11840 ( .B1(n13386), .B2(n13285), .A(n2239), .ZN(n7282) );
  OAI21_X2 U11841 ( .B1(n13457), .B2(n13355), .A(n1747), .ZN(n7315) );
  OAI21_X2 U11842 ( .B1(n13454), .B2(n13356), .A(n1748), .ZN(n7316) );
  OAI21_X2 U11843 ( .B1(n13448), .B2(n13356), .A(n1750), .ZN(n7317) );
  OAI21_X2 U11844 ( .B1(n13445), .B2(n13356), .A(n1751), .ZN(n7318) );
  OAI21_X2 U11845 ( .B1(n13442), .B2(n13356), .A(n1752), .ZN(n7319) );
  OAI21_X2 U11846 ( .B1(n13439), .B2(n13356), .A(n1753), .ZN(n7320) );
  OAI21_X2 U11847 ( .B1(n13436), .B2(n13356), .A(n1754), .ZN(n7321) );
  OAI21_X2 U11848 ( .B1(n13433), .B2(n13356), .A(n1755), .ZN(n7322) );
  OAI21_X2 U11849 ( .B1(n13430), .B2(n13357), .A(n1756), .ZN(n7323) );
  OAI21_X2 U11850 ( .B1(n13427), .B2(n13357), .A(n1757), .ZN(n7324) );
  OAI21_X2 U11851 ( .B1(n13424), .B2(n13356), .A(n1758), .ZN(n7325) );
  OAI21_X2 U11852 ( .B1(n13421), .B2(n13357), .A(n1759), .ZN(n7326) );
  OAI21_X2 U11853 ( .B1(n13415), .B2(n13357), .A(n1761), .ZN(n7327) );
  OAI21_X2 U11854 ( .B1(n13412), .B2(n13357), .A(n1762), .ZN(n7328) );
  OAI21_X2 U11855 ( .B1(n13409), .B2(n13357), .A(n1763), .ZN(n7329) );
  OAI21_X2 U11856 ( .B1(n13406), .B2(n13357), .A(n1764), .ZN(n7330) );
  OAI21_X2 U11857 ( .B1(n13403), .B2(n13356), .A(n1765), .ZN(n7331) );
  OAI21_X2 U11858 ( .B1(n13400), .B2(n13356), .A(n1766), .ZN(n7332) );
  OAI21_X2 U11859 ( .B1(n13397), .B2(n13356), .A(n1767), .ZN(n7333) );
  OAI21_X2 U11860 ( .B1(n13394), .B2(n13355), .A(n1768), .ZN(n7334) );
  OAI21_X2 U11861 ( .B1(n13391), .B2(n13355), .A(n1769), .ZN(n7335) );
  OAI21_X2 U11862 ( .B1(n13388), .B2(n13355), .A(n1770), .ZN(n7336) );
  OAI21_X2 U11863 ( .B1(n13483), .B2(n13355), .A(n1740), .ZN(n7337) );
  OAI21_X2 U11864 ( .B1(n13475), .B2(n13355), .A(n1741), .ZN(n7338) );
  OAI21_X2 U11865 ( .B1(n13472), .B2(n13355), .A(n1742), .ZN(n7339) );
  OAI21_X2 U11866 ( .B1(n13469), .B2(n13355), .A(n1743), .ZN(n7340) );
  OAI21_X2 U11867 ( .B1(n13466), .B2(n13355), .A(n1744), .ZN(n7341) );
  OAI21_X2 U11868 ( .B1(n13463), .B2(n13355), .A(n1745), .ZN(n7342) );
  OAI21_X2 U11869 ( .B1(n13460), .B2(n13355), .A(n1746), .ZN(n7343) );
  OAI21_X2 U11870 ( .B1(n13451), .B2(n13356), .A(n1749), .ZN(n7344) );
  OAI21_X2 U11871 ( .B1(n13418), .B2(n13357), .A(n1760), .ZN(n7345) );
  OAI21_X2 U11872 ( .B1(n13385), .B2(n13355), .A(n1771), .ZN(n7346) );
  OAI21_X2 U11873 ( .B1(n13457), .B2(n13365), .A(n1680), .ZN(n7379) );
  OAI21_X2 U11874 ( .B1(n13454), .B2(n13366), .A(n1681), .ZN(n7380) );
  OAI21_X2 U11875 ( .B1(n13448), .B2(n13366), .A(n1683), .ZN(n7381) );
  OAI21_X2 U11876 ( .B1(n13445), .B2(n13366), .A(n1684), .ZN(n7382) );
  OAI21_X2 U11877 ( .B1(n13442), .B2(n13366), .A(n1685), .ZN(n7383) );
  OAI21_X2 U11878 ( .B1(n13439), .B2(n13366), .A(n1686), .ZN(n7384) );
  OAI21_X2 U11879 ( .B1(n13436), .B2(n13366), .A(n1687), .ZN(n7385) );
  OAI21_X2 U11880 ( .B1(n13433), .B2(n13366), .A(n1688), .ZN(n7386) );
  OAI21_X2 U11881 ( .B1(n13430), .B2(n13367), .A(n1689), .ZN(n7387) );
  OAI21_X2 U11882 ( .B1(n13427), .B2(n13367), .A(n1690), .ZN(n7388) );
  OAI21_X2 U11883 ( .B1(n13424), .B2(n13366), .A(n1691), .ZN(n7389) );
  OAI21_X2 U11884 ( .B1(n13421), .B2(n13367), .A(n1692), .ZN(n7390) );
  OAI21_X2 U11885 ( .B1(n13415), .B2(n13367), .A(n1694), .ZN(n7391) );
  OAI21_X2 U11886 ( .B1(n13412), .B2(n13367), .A(n1695), .ZN(n7392) );
  OAI21_X2 U11887 ( .B1(n13409), .B2(n13367), .A(n1696), .ZN(n7393) );
  OAI21_X2 U11888 ( .B1(n13406), .B2(n13367), .A(n1697), .ZN(n7394) );
  OAI21_X2 U11889 ( .B1(n13403), .B2(n13366), .A(n1698), .ZN(n7395) );
  OAI21_X2 U11890 ( .B1(n13400), .B2(n13366), .A(n1699), .ZN(n7396) );
  OAI21_X2 U11891 ( .B1(n13397), .B2(n13366), .A(n1700), .ZN(n7397) );
  OAI21_X2 U11892 ( .B1(n13394), .B2(n13365), .A(n1701), .ZN(n7398) );
  OAI21_X2 U11893 ( .B1(n13391), .B2(n13365), .A(n1702), .ZN(n7399) );
  OAI21_X2 U11894 ( .B1(n13388), .B2(n13365), .A(n1703), .ZN(n7400) );
  OAI21_X2 U11895 ( .B1(n13483), .B2(n13365), .A(n1673), .ZN(n7401) );
  OAI21_X2 U11896 ( .B1(n13475), .B2(n13365), .A(n1674), .ZN(n7402) );
  OAI21_X2 U11897 ( .B1(n13472), .B2(n13365), .A(n1675), .ZN(n7403) );
  OAI21_X2 U11898 ( .B1(n13469), .B2(n13365), .A(n1676), .ZN(n7404) );
  OAI21_X2 U11899 ( .B1(n13466), .B2(n13365), .A(n1677), .ZN(n7405) );
  OAI21_X2 U11900 ( .B1(n13463), .B2(n13365), .A(n1678), .ZN(n7406) );
  OAI21_X2 U11901 ( .B1(n13460), .B2(n13365), .A(n1679), .ZN(n7407) );
  OAI21_X2 U11902 ( .B1(n13451), .B2(n13366), .A(n1682), .ZN(n7408) );
  OAI21_X2 U11903 ( .B1(n13418), .B2(n13367), .A(n1693), .ZN(n7409) );
  OAI21_X2 U11904 ( .B1(n13385), .B2(n13365), .A(n1704), .ZN(n7410) );
  OAI21_X2 U11905 ( .B1(n13457), .B2(n13375), .A(n1613), .ZN(n7443) );
  OAI21_X2 U11906 ( .B1(n13454), .B2(n13376), .A(n1614), .ZN(n7444) );
  OAI21_X2 U11907 ( .B1(n13448), .B2(n13376), .A(n1616), .ZN(n7445) );
  OAI21_X2 U11908 ( .B1(n13445), .B2(n13376), .A(n1617), .ZN(n7446) );
  OAI21_X2 U11909 ( .B1(n13442), .B2(n13376), .A(n1618), .ZN(n7447) );
  OAI21_X2 U11910 ( .B1(n13439), .B2(n13376), .A(n1619), .ZN(n7448) );
  OAI21_X2 U11911 ( .B1(n13436), .B2(n13376), .A(n1620), .ZN(n7449) );
  OAI21_X2 U11912 ( .B1(n13433), .B2(n13376), .A(n1621), .ZN(n7450) );
  OAI21_X2 U11913 ( .B1(n13430), .B2(n13377), .A(n1622), .ZN(n7451) );
  OAI21_X2 U11914 ( .B1(n13427), .B2(n13377), .A(n1623), .ZN(n7452) );
  OAI21_X2 U11915 ( .B1(n13424), .B2(n13376), .A(n1624), .ZN(n7453) );
  OAI21_X2 U11916 ( .B1(n13421), .B2(n13377), .A(n1625), .ZN(n7454) );
  OAI21_X2 U11917 ( .B1(n13415), .B2(n13377), .A(n1627), .ZN(n7455) );
  OAI21_X2 U11918 ( .B1(n13412), .B2(n13377), .A(n1628), .ZN(n7456) );
  OAI21_X2 U11919 ( .B1(n13409), .B2(n13377), .A(n1629), .ZN(n7457) );
  OAI21_X2 U11920 ( .B1(n13406), .B2(n13377), .A(n1630), .ZN(n7458) );
  OAI21_X2 U11921 ( .B1(n13403), .B2(n13376), .A(n1631), .ZN(n7459) );
  OAI21_X2 U11922 ( .B1(n13400), .B2(n13376), .A(n1632), .ZN(n7460) );
  OAI21_X2 U11923 ( .B1(n13397), .B2(n13376), .A(n1633), .ZN(n7461) );
  OAI21_X2 U11924 ( .B1(n13394), .B2(n13375), .A(n1634), .ZN(n7462) );
  OAI21_X2 U11925 ( .B1(n13391), .B2(n13375), .A(n1635), .ZN(n7463) );
  OAI21_X2 U11926 ( .B1(n13388), .B2(n13375), .A(n1636), .ZN(n7464) );
  OAI21_X2 U11927 ( .B1(n13483), .B2(n13375), .A(n1606), .ZN(n7465) );
  OAI21_X2 U11928 ( .B1(n13475), .B2(n13375), .A(n1607), .ZN(n7466) );
  OAI21_X2 U11929 ( .B1(n13472), .B2(n13375), .A(n1608), .ZN(n7467) );
  OAI21_X2 U11930 ( .B1(n13469), .B2(n13375), .A(n1609), .ZN(n7468) );
  OAI21_X2 U11931 ( .B1(n13466), .B2(n13375), .A(n1610), .ZN(n7469) );
  OAI21_X2 U11932 ( .B1(n13463), .B2(n13375), .A(n1611), .ZN(n7470) );
  OAI21_X2 U11933 ( .B1(n13460), .B2(n13375), .A(n1612), .ZN(n7471) );
  OAI21_X2 U11934 ( .B1(n13451), .B2(n13376), .A(n1615), .ZN(n7472) );
  OAI21_X2 U11935 ( .B1(n13418), .B2(n13377), .A(n1626), .ZN(n7473) );
  OAI21_X2 U11936 ( .B1(n13385), .B2(n13375), .A(n1637), .ZN(n7474) );
  OAI21_X2 U11937 ( .B1(n13457), .B2(n13478), .A(n1522), .ZN(n7507) );
  OAI21_X2 U11938 ( .B1(n13454), .B2(n13479), .A(n1524), .ZN(n7508) );
  OAI21_X2 U11939 ( .B1(n13448), .B2(n13479), .A(n1528), .ZN(n7509) );
  OAI21_X2 U11940 ( .B1(n13445), .B2(n13479), .A(n1530), .ZN(n7510) );
  OAI21_X2 U11941 ( .B1(n13442), .B2(n13479), .A(n1532), .ZN(n7511) );
  OAI21_X2 U11942 ( .B1(n13439), .B2(n13479), .A(n1534), .ZN(n7512) );
  OAI21_X2 U11943 ( .B1(n13436), .B2(n13479), .A(n1536), .ZN(n7513) );
  OAI21_X2 U11944 ( .B1(n13433), .B2(n13479), .A(n1538), .ZN(n7514) );
  OAI21_X2 U11945 ( .B1(n13430), .B2(n13480), .A(n1540), .ZN(n7515) );
  OAI21_X2 U11946 ( .B1(n13427), .B2(n13480), .A(n1542), .ZN(n7516) );
  OAI21_X2 U11947 ( .B1(n13424), .B2(n13479), .A(n1544), .ZN(n7517) );
  OAI21_X2 U11948 ( .B1(n13421), .B2(n13480), .A(n1546), .ZN(n7518) );
  OAI21_X2 U11949 ( .B1(n13415), .B2(n13480), .A(n1550), .ZN(n7519) );
  OAI21_X2 U11950 ( .B1(n13412), .B2(n13480), .A(n1552), .ZN(n7520) );
  OAI21_X2 U11951 ( .B1(n13409), .B2(n13480), .A(n1554), .ZN(n7521) );
  OAI21_X2 U11952 ( .B1(n13406), .B2(n13480), .A(n1556), .ZN(n7522) );
  OAI21_X2 U11953 ( .B1(n13403), .B2(n13479), .A(n1558), .ZN(n7523) );
  OAI21_X2 U11954 ( .B1(n13400), .B2(n13479), .A(n1560), .ZN(n7524) );
  OAI21_X2 U11955 ( .B1(n13397), .B2(n13479), .A(n1562), .ZN(n7525) );
  OAI21_X2 U11956 ( .B1(n13394), .B2(n13478), .A(n1564), .ZN(n7526) );
  OAI21_X2 U11957 ( .B1(n13391), .B2(n13478), .A(n1566), .ZN(n7527) );
  OAI21_X2 U11958 ( .B1(n13388), .B2(n13478), .A(n1568), .ZN(n7528) );
  OAI21_X2 U11959 ( .B1(n13483), .B2(n13478), .A(n1508), .ZN(n7529) );
  OAI21_X2 U11960 ( .B1(n13475), .B2(n13478), .A(n1510), .ZN(n7530) );
  OAI21_X2 U11961 ( .B1(n13472), .B2(n13478), .A(n1512), .ZN(n7531) );
  OAI21_X2 U11962 ( .B1(n13469), .B2(n13478), .A(n1514), .ZN(n7532) );
  OAI21_X2 U11963 ( .B1(n13466), .B2(n13478), .A(n1516), .ZN(n7533) );
  OAI21_X2 U11964 ( .B1(n13463), .B2(n13478), .A(n1518), .ZN(n7534) );
  OAI21_X2 U11965 ( .B1(n13460), .B2(n13478), .A(n1520), .ZN(n7535) );
  OAI21_X2 U11966 ( .B1(n13451), .B2(n13479), .A(n1526), .ZN(n7536) );
  OAI21_X2 U11967 ( .B1(n13418), .B2(n13480), .A(n1548), .ZN(n7537) );
  OAI21_X2 U11968 ( .B1(n13385), .B2(n13478), .A(n1570), .ZN(n7538) );
  OAI21_X2 U11969 ( .B1(n1521), .B2(n13240), .A(n2517), .ZN(n7571) );
  OAI21_X2 U11970 ( .B1(n1523), .B2(n13241), .A(n2518), .ZN(n7572) );
  OAI21_X2 U11971 ( .B1(n1527), .B2(n13241), .A(n2520), .ZN(n7573) );
  OAI21_X2 U11972 ( .B1(n1529), .B2(n13241), .A(n2521), .ZN(n7574) );
  OAI21_X2 U11973 ( .B1(n1531), .B2(n13241), .A(n2522), .ZN(n7575) );
  OAI21_X2 U11974 ( .B1(n1533), .B2(n13241), .A(n2523), .ZN(n7576) );
  OAI21_X2 U11975 ( .B1(n1535), .B2(n13241), .A(n2524), .ZN(n7577) );
  OAI21_X2 U11976 ( .B1(n1537), .B2(n13241), .A(n2525), .ZN(n7578) );
  OAI21_X2 U11977 ( .B1(n1539), .B2(n13242), .A(n2526), .ZN(n7579) );
  OAI21_X2 U11978 ( .B1(n1541), .B2(n13242), .A(n2527), .ZN(n7580) );
  OAI21_X2 U11979 ( .B1(n1543), .B2(n13241), .A(n2528), .ZN(n7581) );
  OAI21_X2 U11980 ( .B1(n1545), .B2(n13242), .A(n2529), .ZN(n7582) );
  OAI21_X2 U11981 ( .B1(n1549), .B2(n13242), .A(n2531), .ZN(n7583) );
  OAI21_X2 U11982 ( .B1(n1551), .B2(n13242), .A(n2532), .ZN(n7584) );
  OAI21_X2 U11983 ( .B1(n1553), .B2(n13242), .A(n2533), .ZN(n7585) );
  OAI21_X2 U11984 ( .B1(n1555), .B2(n13242), .A(n2534), .ZN(n7586) );
  OAI21_X2 U11985 ( .B1(n1557), .B2(n13241), .A(n2535), .ZN(n7587) );
  OAI21_X2 U11986 ( .B1(n1559), .B2(n13241), .A(n2536), .ZN(n7588) );
  OAI21_X2 U11987 ( .B1(n1561), .B2(n13241), .A(n2537), .ZN(n7589) );
  OAI21_X2 U11988 ( .B1(n1563), .B2(n13240), .A(n2538), .ZN(n7590) );
  OAI21_X2 U11989 ( .B1(n1565), .B2(n13240), .A(n2539), .ZN(n7591) );
  OAI21_X2 U11990 ( .B1(n1567), .B2(n13240), .A(n2540), .ZN(n7592) );
  OAI21_X2 U11991 ( .B1(n1506), .B2(n13240), .A(n2510), .ZN(n7593) );
  OAI21_X2 U11992 ( .B1(n1509), .B2(n13240), .A(n2511), .ZN(n7594) );
  OAI21_X2 U11993 ( .B1(n1511), .B2(n13240), .A(n2512), .ZN(n7595) );
  OAI21_X2 U11994 ( .B1(n1513), .B2(n13240), .A(n2513), .ZN(n7596) );
  OAI21_X2 U11995 ( .B1(n1515), .B2(n13240), .A(n2514), .ZN(n7597) );
  OAI21_X2 U11996 ( .B1(n1517), .B2(n13240), .A(n2515), .ZN(n7598) );
  OAI21_X2 U11997 ( .B1(n1519), .B2(n13240), .A(n2516), .ZN(n7599) );
  OAI21_X2 U11998 ( .B1(n1525), .B2(n13241), .A(n2519), .ZN(n7600) );
  OAI21_X2 U11999 ( .B1(n1547), .B2(n13242), .A(n2530), .ZN(n7601) );
  OAI21_X2 U12000 ( .B1(n1569), .B2(n13240), .A(n2541), .ZN(n7602) );
  OAI21_X2 U12001 ( .B1(n1521), .B2(n13250), .A(n2449), .ZN(n7635) );
  OAI21_X2 U12002 ( .B1(n1523), .B2(n13251), .A(n2450), .ZN(n7636) );
  OAI21_X2 U12003 ( .B1(n1527), .B2(n13251), .A(n2452), .ZN(n7637) );
  OAI21_X2 U12004 ( .B1(n1529), .B2(n13251), .A(n2453), .ZN(n7638) );
  OAI21_X2 U12005 ( .B1(n1531), .B2(n13251), .A(n2454), .ZN(n7639) );
  OAI21_X2 U12006 ( .B1(n1533), .B2(n13251), .A(n2455), .ZN(n7640) );
  OAI21_X2 U12007 ( .B1(n1535), .B2(n13251), .A(n2456), .ZN(n7641) );
  OAI21_X2 U12008 ( .B1(n1537), .B2(n13251), .A(n2457), .ZN(n7642) );
  OAI21_X2 U12009 ( .B1(n1539), .B2(n13252), .A(n2458), .ZN(n7643) );
  OAI21_X2 U12010 ( .B1(n1541), .B2(n13252), .A(n2459), .ZN(n7644) );
  OAI21_X2 U12011 ( .B1(n1543), .B2(n13251), .A(n2460), .ZN(n7645) );
  OAI21_X2 U12012 ( .B1(n1545), .B2(n13252), .A(n2461), .ZN(n7646) );
  OAI21_X2 U12013 ( .B1(n1549), .B2(n13252), .A(n2463), .ZN(n7647) );
  OAI21_X2 U12014 ( .B1(n1551), .B2(n13252), .A(n2464), .ZN(n7648) );
  OAI21_X2 U12015 ( .B1(n1553), .B2(n13252), .A(n2465), .ZN(n7649) );
  OAI21_X2 U12016 ( .B1(n1555), .B2(n13252), .A(n2466), .ZN(n7650) );
  OAI21_X2 U12017 ( .B1(n1557), .B2(n13251), .A(n2467), .ZN(n7651) );
  OAI21_X2 U12018 ( .B1(n1559), .B2(n13251), .A(n2468), .ZN(n7652) );
  OAI21_X2 U12019 ( .B1(n1561), .B2(n13251), .A(n2469), .ZN(n7653) );
  OAI21_X2 U12020 ( .B1(n1563), .B2(n13250), .A(n2470), .ZN(n7654) );
  OAI21_X2 U12021 ( .B1(n1565), .B2(n13250), .A(n2471), .ZN(n7655) );
  OAI21_X2 U12022 ( .B1(n1567), .B2(n13250), .A(n2472), .ZN(n7656) );
  OAI21_X2 U12023 ( .B1(n1506), .B2(n13250), .A(n2442), .ZN(n7657) );
  OAI21_X2 U12024 ( .B1(n1509), .B2(n13250), .A(n2443), .ZN(n7658) );
  OAI21_X2 U12025 ( .B1(n1511), .B2(n13250), .A(n2444), .ZN(n7659) );
  OAI21_X2 U12026 ( .B1(n1513), .B2(n13250), .A(n2445), .ZN(n7660) );
  OAI21_X2 U12027 ( .B1(n1515), .B2(n13250), .A(n2446), .ZN(n7661) );
  OAI21_X2 U12028 ( .B1(n1517), .B2(n13250), .A(n2447), .ZN(n7662) );
  OAI21_X2 U12029 ( .B1(n1519), .B2(n13250), .A(n2448), .ZN(n7663) );
  OAI21_X2 U12030 ( .B1(n1525), .B2(n13251), .A(n2451), .ZN(n7664) );
  OAI21_X2 U12031 ( .B1(n1547), .B2(n13252), .A(n2462), .ZN(n7665) );
  OAI21_X2 U12032 ( .B1(n1569), .B2(n13250), .A(n2473), .ZN(n7666) );
  OAI21_X2 U12033 ( .B1(n1521), .B2(n13260), .A(n2382), .ZN(n7699) );
  OAI21_X2 U12034 ( .B1(n1523), .B2(n13261), .A(n2383), .ZN(n7700) );
  OAI21_X2 U12035 ( .B1(n1527), .B2(n13261), .A(n2385), .ZN(n7701) );
  OAI21_X2 U12036 ( .B1(n1529), .B2(n13261), .A(n2386), .ZN(n7702) );
  OAI21_X2 U12037 ( .B1(n1531), .B2(n13261), .A(n2387), .ZN(n7703) );
  OAI21_X2 U12038 ( .B1(n1533), .B2(n13261), .A(n2388), .ZN(n7704) );
  OAI21_X2 U12039 ( .B1(n1535), .B2(n13261), .A(n2389), .ZN(n7705) );
  OAI21_X2 U12040 ( .B1(n1537), .B2(n13261), .A(n2390), .ZN(n7706) );
  OAI21_X2 U12041 ( .B1(n1539), .B2(n13262), .A(n2391), .ZN(n7707) );
  OAI21_X2 U12042 ( .B1(n1541), .B2(n13262), .A(n2392), .ZN(n7708) );
  OAI21_X2 U12043 ( .B1(n1543), .B2(n13261), .A(n2393), .ZN(n7709) );
  OAI21_X2 U12044 ( .B1(n1545), .B2(n13262), .A(n2394), .ZN(n7710) );
  OAI21_X2 U12045 ( .B1(n1549), .B2(n13262), .A(n2396), .ZN(n7711) );
  OAI21_X2 U12046 ( .B1(n1551), .B2(n13262), .A(n2397), .ZN(n7712) );
  OAI21_X2 U12047 ( .B1(n1553), .B2(n13262), .A(n2398), .ZN(n7713) );
  OAI21_X2 U12048 ( .B1(n1555), .B2(n13262), .A(n2399), .ZN(n7714) );
  OAI21_X2 U12049 ( .B1(n1557), .B2(n13261), .A(n2400), .ZN(n7715) );
  OAI21_X2 U12050 ( .B1(n1559), .B2(n13261), .A(n2401), .ZN(n7716) );
  OAI21_X2 U12051 ( .B1(n1561), .B2(n13261), .A(n2402), .ZN(n7717) );
  OAI21_X2 U12052 ( .B1(n1563), .B2(n13260), .A(n2403), .ZN(n7718) );
  OAI21_X2 U12053 ( .B1(n1565), .B2(n13260), .A(n2404), .ZN(n7719) );
  OAI21_X2 U12054 ( .B1(n1567), .B2(n13260), .A(n2405), .ZN(n7720) );
  OAI21_X2 U12055 ( .B1(n1506), .B2(n13260), .A(n2375), .ZN(n7721) );
  OAI21_X2 U12056 ( .B1(n1509), .B2(n13260), .A(n2376), .ZN(n7722) );
  OAI21_X2 U12057 ( .B1(n1511), .B2(n13260), .A(n2377), .ZN(n7723) );
  OAI21_X2 U12058 ( .B1(n1513), .B2(n13260), .A(n2378), .ZN(n7724) );
  OAI21_X2 U12059 ( .B1(n1515), .B2(n13260), .A(n2379), .ZN(n7725) );
  OAI21_X2 U12060 ( .B1(n1517), .B2(n13260), .A(n2380), .ZN(n7726) );
  OAI21_X2 U12061 ( .B1(n1519), .B2(n13260), .A(n2381), .ZN(n7727) );
  OAI21_X2 U12062 ( .B1(n1525), .B2(n13261), .A(n2384), .ZN(n7728) );
  OAI21_X2 U12063 ( .B1(n1547), .B2(n13262), .A(n2395), .ZN(n7729) );
  OAI21_X2 U12064 ( .B1(n1569), .B2(n13260), .A(n2406), .ZN(n7730) );
  OAI21_X2 U12065 ( .B1(n13458), .B2(n13270), .A(n2315), .ZN(n7763) );
  OAI21_X2 U12066 ( .B1(n13455), .B2(n13271), .A(n2316), .ZN(n7764) );
  OAI21_X2 U12067 ( .B1(n13449), .B2(n13271), .A(n2318), .ZN(n7765) );
  OAI21_X2 U12068 ( .B1(n13446), .B2(n13271), .A(n2319), .ZN(n7766) );
  OAI21_X2 U12069 ( .B1(n13443), .B2(n13271), .A(n2320), .ZN(n7767) );
  OAI21_X2 U12070 ( .B1(n13440), .B2(n13271), .A(n2321), .ZN(n7768) );
  OAI21_X2 U12071 ( .B1(n13437), .B2(n13271), .A(n2322), .ZN(n7769) );
  OAI21_X2 U12072 ( .B1(n13434), .B2(n13271), .A(n2323), .ZN(n7770) );
  OAI21_X2 U12073 ( .B1(n13431), .B2(n13272), .A(n2324), .ZN(n7771) );
  OAI21_X2 U12074 ( .B1(n13428), .B2(n13272), .A(n2325), .ZN(n7772) );
  OAI21_X2 U12075 ( .B1(n13425), .B2(n13271), .A(n2326), .ZN(n7773) );
  OAI21_X2 U12076 ( .B1(n13422), .B2(n13272), .A(n2327), .ZN(n7774) );
  OAI21_X2 U12077 ( .B1(n13416), .B2(n13272), .A(n2329), .ZN(n7775) );
  OAI21_X2 U12078 ( .B1(n13413), .B2(n13272), .A(n2330), .ZN(n7776) );
  OAI21_X2 U12079 ( .B1(n13410), .B2(n13272), .A(n2331), .ZN(n7777) );
  OAI21_X2 U12080 ( .B1(n13407), .B2(n13272), .A(n2332), .ZN(n7778) );
  OAI21_X2 U12081 ( .B1(n13404), .B2(n13271), .A(n2333), .ZN(n7779) );
  OAI21_X2 U12082 ( .B1(n13401), .B2(n13271), .A(n2334), .ZN(n7780) );
  OAI21_X2 U12083 ( .B1(n13398), .B2(n13271), .A(n2335), .ZN(n7781) );
  OAI21_X2 U12084 ( .B1(n13395), .B2(n13270), .A(n2336), .ZN(n7782) );
  OAI21_X2 U12085 ( .B1(n13392), .B2(n13270), .A(n2337), .ZN(n7783) );
  OAI21_X2 U12086 ( .B1(n13389), .B2(n13270), .A(n2338), .ZN(n7784) );
  OAI21_X2 U12087 ( .B1(n13484), .B2(n13270), .A(n2308), .ZN(n7785) );
  OAI21_X2 U12088 ( .B1(n13476), .B2(n13270), .A(n2309), .ZN(n7786) );
  OAI21_X2 U12089 ( .B1(n13473), .B2(n13270), .A(n2310), .ZN(n7787) );
  OAI21_X2 U12090 ( .B1(n13470), .B2(n13270), .A(n2311), .ZN(n7788) );
  OAI21_X2 U12091 ( .B1(n13467), .B2(n13270), .A(n2312), .ZN(n7789) );
  OAI21_X2 U12092 ( .B1(n13464), .B2(n13270), .A(n2313), .ZN(n7790) );
  OAI21_X2 U12093 ( .B1(n13461), .B2(n13270), .A(n2314), .ZN(n7791) );
  OAI21_X2 U12094 ( .B1(n13452), .B2(n13271), .A(n2317), .ZN(n7792) );
  OAI21_X2 U12095 ( .B1(n13419), .B2(n13272), .A(n2328), .ZN(n7793) );
  OAI21_X2 U12096 ( .B1(n13386), .B2(n13270), .A(n2339), .ZN(n7794) );
  OAI21_X2 U12097 ( .B1(n13458), .B2(n13280), .A(n2248), .ZN(n7827) );
  OAI21_X2 U12098 ( .B1(n13455), .B2(n13281), .A(n2249), .ZN(n7828) );
  OAI21_X2 U12099 ( .B1(n13449), .B2(n13281), .A(n2251), .ZN(n7829) );
  OAI21_X2 U12100 ( .B1(n13446), .B2(n13281), .A(n2252), .ZN(n7830) );
  OAI21_X2 U12101 ( .B1(n13443), .B2(n13281), .A(n2253), .ZN(n7831) );
  OAI21_X2 U12102 ( .B1(n13440), .B2(n13281), .A(n2254), .ZN(n7832) );
  OAI21_X2 U12103 ( .B1(n13437), .B2(n13281), .A(n2255), .ZN(n7833) );
  OAI21_X2 U12104 ( .B1(n13434), .B2(n13281), .A(n2256), .ZN(n7834) );
  OAI21_X2 U12105 ( .B1(n13431), .B2(n13282), .A(n2257), .ZN(n7835) );
  OAI21_X2 U12106 ( .B1(n13428), .B2(n13282), .A(n2258), .ZN(n7836) );
  OAI21_X2 U12107 ( .B1(n13425), .B2(n13281), .A(n2259), .ZN(n7837) );
  OAI21_X2 U12108 ( .B1(n13422), .B2(n13282), .A(n2260), .ZN(n7838) );
  OAI21_X2 U12109 ( .B1(n13416), .B2(n13282), .A(n2262), .ZN(n7839) );
  OAI21_X2 U12110 ( .B1(n13413), .B2(n13282), .A(n2263), .ZN(n7840) );
  OAI21_X2 U12111 ( .B1(n13410), .B2(n13282), .A(n2264), .ZN(n7841) );
  OAI21_X2 U12112 ( .B1(n13407), .B2(n13282), .A(n2265), .ZN(n7842) );
  OAI21_X2 U12113 ( .B1(n13404), .B2(n13281), .A(n2266), .ZN(n7843) );
  OAI21_X2 U12114 ( .B1(n13401), .B2(n13281), .A(n2267), .ZN(n7844) );
  OAI21_X2 U12115 ( .B1(n13398), .B2(n13281), .A(n2268), .ZN(n7845) );
  OAI21_X2 U12116 ( .B1(n13395), .B2(n13280), .A(n2269), .ZN(n7846) );
  OAI21_X2 U12117 ( .B1(n13392), .B2(n13280), .A(n2270), .ZN(n7847) );
  OAI21_X2 U12118 ( .B1(n13389), .B2(n13280), .A(n2271), .ZN(n7848) );
  OAI21_X2 U12119 ( .B1(n13484), .B2(n13280), .A(n2241), .ZN(n7849) );
  OAI21_X2 U12120 ( .B1(n13476), .B2(n13280), .A(n2242), .ZN(n7850) );
  OAI21_X2 U12121 ( .B1(n13473), .B2(n13280), .A(n2243), .ZN(n7851) );
  OAI21_X2 U12122 ( .B1(n13470), .B2(n13280), .A(n2244), .ZN(n7852) );
  OAI21_X2 U12123 ( .B1(n13467), .B2(n13280), .A(n2245), .ZN(n7853) );
  OAI21_X2 U12124 ( .B1(n13464), .B2(n13280), .A(n2246), .ZN(n7854) );
  OAI21_X2 U12125 ( .B1(n13461), .B2(n13280), .A(n2247), .ZN(n7855) );
  OAI21_X2 U12126 ( .B1(n13452), .B2(n13281), .A(n2250), .ZN(n7856) );
  OAI21_X2 U12127 ( .B1(n13419), .B2(n13282), .A(n2261), .ZN(n7857) );
  OAI21_X2 U12128 ( .B1(n13386), .B2(n13280), .A(n2272), .ZN(n7858) );
  OAI21_X2 U12129 ( .B1(n13458), .B2(n13295), .A(n2148), .ZN(n7891) );
  OAI21_X2 U12130 ( .B1(n13455), .B2(n13296), .A(n2149), .ZN(n7892) );
  OAI21_X2 U12131 ( .B1(n13449), .B2(n13296), .A(n2151), .ZN(n7893) );
  OAI21_X2 U12132 ( .B1(n13446), .B2(n13296), .A(n2152), .ZN(n7894) );
  OAI21_X2 U12133 ( .B1(n13443), .B2(n13296), .A(n2153), .ZN(n7895) );
  OAI21_X2 U12134 ( .B1(n13440), .B2(n13296), .A(n2154), .ZN(n7896) );
  OAI21_X2 U12135 ( .B1(n13437), .B2(n13296), .A(n2155), .ZN(n7897) );
  OAI21_X2 U12136 ( .B1(n13434), .B2(n13296), .A(n2156), .ZN(n7898) );
  OAI21_X2 U12137 ( .B1(n13431), .B2(n13297), .A(n2157), .ZN(n7899) );
  OAI21_X2 U12138 ( .B1(n13428), .B2(n13297), .A(n2158), .ZN(n7900) );
  OAI21_X2 U12139 ( .B1(n13425), .B2(n13296), .A(n2159), .ZN(n7901) );
  OAI21_X2 U12140 ( .B1(n13422), .B2(n13297), .A(n2160), .ZN(n7902) );
  OAI21_X2 U12141 ( .B1(n13416), .B2(n13297), .A(n2162), .ZN(n7903) );
  OAI21_X2 U12142 ( .B1(n13413), .B2(n13297), .A(n2163), .ZN(n7904) );
  OAI21_X2 U12143 ( .B1(n13410), .B2(n13297), .A(n2164), .ZN(n7905) );
  OAI21_X2 U12144 ( .B1(n13407), .B2(n13297), .A(n2165), .ZN(n7906) );
  OAI21_X2 U12145 ( .B1(n13404), .B2(n13296), .A(n2166), .ZN(n7907) );
  OAI21_X2 U12146 ( .B1(n13401), .B2(n13296), .A(n2167), .ZN(n7908) );
  OAI21_X2 U12147 ( .B1(n13398), .B2(n13296), .A(n2168), .ZN(n7909) );
  OAI21_X2 U12148 ( .B1(n13395), .B2(n13295), .A(n2169), .ZN(n7910) );
  OAI21_X2 U12149 ( .B1(n13392), .B2(n13295), .A(n2170), .ZN(n7911) );
  OAI21_X2 U12150 ( .B1(n13389), .B2(n13295), .A(n2171), .ZN(n7912) );
  OAI21_X2 U12151 ( .B1(n13484), .B2(n13295), .A(n2141), .ZN(n7913) );
  OAI21_X2 U12152 ( .B1(n13476), .B2(n13295), .A(n2142), .ZN(n7914) );
  OAI21_X2 U12153 ( .B1(n13473), .B2(n13295), .A(n2143), .ZN(n7915) );
  OAI21_X2 U12154 ( .B1(n13470), .B2(n13295), .A(n2144), .ZN(n7916) );
  OAI21_X2 U12155 ( .B1(n13467), .B2(n13295), .A(n2145), .ZN(n7917) );
  OAI21_X2 U12156 ( .B1(n13464), .B2(n13295), .A(n2146), .ZN(n7918) );
  OAI21_X2 U12157 ( .B1(n13461), .B2(n13295), .A(n2147), .ZN(n7919) );
  OAI21_X2 U12158 ( .B1(n13452), .B2(n13296), .A(n2150), .ZN(n7920) );
  OAI21_X2 U12159 ( .B1(n13419), .B2(n13297), .A(n2161), .ZN(n7921) );
  OAI21_X2 U12160 ( .B1(n13386), .B2(n13295), .A(n2172), .ZN(n7922) );
  OAI21_X2 U12161 ( .B1(n13458), .B2(n13305), .A(n2081), .ZN(n7955) );
  OAI21_X2 U12162 ( .B1(n13455), .B2(n13306), .A(n2082), .ZN(n7956) );
  OAI21_X2 U12163 ( .B1(n13449), .B2(n13306), .A(n2084), .ZN(n7957) );
  OAI21_X2 U12164 ( .B1(n13446), .B2(n13306), .A(n2085), .ZN(n7958) );
  OAI21_X2 U12165 ( .B1(n13443), .B2(n13306), .A(n2086), .ZN(n7959) );
  OAI21_X2 U12166 ( .B1(n13440), .B2(n13306), .A(n2087), .ZN(n7960) );
  OAI21_X2 U12167 ( .B1(n13437), .B2(n13306), .A(n2088), .ZN(n7961) );
  OAI21_X2 U12168 ( .B1(n13434), .B2(n13306), .A(n2089), .ZN(n7962) );
  OAI21_X2 U12169 ( .B1(n13431), .B2(n13307), .A(n2090), .ZN(n7963) );
  OAI21_X2 U12170 ( .B1(n13428), .B2(n13307), .A(n2091), .ZN(n7964) );
  OAI21_X2 U12171 ( .B1(n13425), .B2(n13306), .A(n2092), .ZN(n7965) );
  OAI21_X2 U12172 ( .B1(n13422), .B2(n13307), .A(n2093), .ZN(n7966) );
  OAI21_X2 U12173 ( .B1(n13416), .B2(n13307), .A(n2095), .ZN(n7967) );
  OAI21_X2 U12174 ( .B1(n13413), .B2(n13307), .A(n2096), .ZN(n7968) );
  OAI21_X2 U12175 ( .B1(n13410), .B2(n13307), .A(n2097), .ZN(n7969) );
  OAI21_X2 U12176 ( .B1(n13407), .B2(n13307), .A(n2098), .ZN(n7970) );
  OAI21_X2 U12177 ( .B1(n13404), .B2(n13306), .A(n2099), .ZN(n7971) );
  OAI21_X2 U12178 ( .B1(n13401), .B2(n13306), .A(n2100), .ZN(n7972) );
  OAI21_X2 U12179 ( .B1(n13398), .B2(n13306), .A(n2101), .ZN(n7973) );
  OAI21_X2 U12180 ( .B1(n13395), .B2(n13305), .A(n2102), .ZN(n7974) );
  OAI21_X2 U12181 ( .B1(n13392), .B2(n13305), .A(n2103), .ZN(n7975) );
  OAI21_X2 U12182 ( .B1(n13389), .B2(n13305), .A(n2104), .ZN(n7976) );
  OAI21_X2 U12183 ( .B1(n13484), .B2(n13305), .A(n2074), .ZN(n7977) );
  OAI21_X2 U12184 ( .B1(n13476), .B2(n13305), .A(n2075), .ZN(n7978) );
  OAI21_X2 U12185 ( .B1(n13473), .B2(n13305), .A(n2076), .ZN(n7979) );
  OAI21_X2 U12186 ( .B1(n13470), .B2(n13305), .A(n2077), .ZN(n7980) );
  OAI21_X2 U12187 ( .B1(n13467), .B2(n13305), .A(n2078), .ZN(n7981) );
  OAI21_X2 U12188 ( .B1(n13464), .B2(n13305), .A(n2079), .ZN(n7982) );
  OAI21_X2 U12189 ( .B1(n13461), .B2(n13305), .A(n2080), .ZN(n7983) );
  OAI21_X2 U12190 ( .B1(n13452), .B2(n13306), .A(n2083), .ZN(n7984) );
  OAI21_X2 U12191 ( .B1(n13419), .B2(n13307), .A(n2094), .ZN(n7985) );
  OAI21_X2 U12192 ( .B1(n13386), .B2(n13305), .A(n2105), .ZN(n7986) );
  OAI21_X2 U12193 ( .B1(n13458), .B2(n13315), .A(n2015), .ZN(n8019) );
  OAI21_X2 U12194 ( .B1(n13455), .B2(n13316), .A(n2016), .ZN(n8020) );
  OAI21_X2 U12195 ( .B1(n13449), .B2(n13316), .A(n2018), .ZN(n8021) );
  OAI21_X2 U12196 ( .B1(n13446), .B2(n13316), .A(n2019), .ZN(n8022) );
  OAI21_X2 U12197 ( .B1(n13443), .B2(n13316), .A(n2020), .ZN(n8023) );
  OAI21_X2 U12198 ( .B1(n13440), .B2(n13316), .A(n2021), .ZN(n8024) );
  OAI21_X2 U12199 ( .B1(n13437), .B2(n13316), .A(n2022), .ZN(n8025) );
  OAI21_X2 U12200 ( .B1(n13434), .B2(n13316), .A(n2023), .ZN(n8026) );
  OAI21_X2 U12201 ( .B1(n13431), .B2(n13317), .A(n2024), .ZN(n8027) );
  OAI21_X2 U12202 ( .B1(n13428), .B2(n13317), .A(n2025), .ZN(n8028) );
  OAI21_X2 U12203 ( .B1(n13425), .B2(n13316), .A(n2026), .ZN(n8029) );
  OAI21_X2 U12204 ( .B1(n13422), .B2(n13317), .A(n2027), .ZN(n8030) );
  OAI21_X2 U12205 ( .B1(n13416), .B2(n13317), .A(n2029), .ZN(n8031) );
  OAI21_X2 U12206 ( .B1(n13413), .B2(n13317), .A(n2030), .ZN(n8032) );
  OAI21_X2 U12207 ( .B1(n13410), .B2(n13317), .A(n2031), .ZN(n8033) );
  OAI21_X2 U12208 ( .B1(n13407), .B2(n13317), .A(n2032), .ZN(n8034) );
  OAI21_X2 U12209 ( .B1(n13404), .B2(n13316), .A(n2033), .ZN(n8035) );
  OAI21_X2 U12210 ( .B1(n13401), .B2(n13316), .A(n2034), .ZN(n8036) );
  OAI21_X2 U12211 ( .B1(n13398), .B2(n13316), .A(n2035), .ZN(n8037) );
  OAI21_X2 U12212 ( .B1(n13395), .B2(n13315), .A(n2036), .ZN(n8038) );
  OAI21_X2 U12213 ( .B1(n13392), .B2(n13315), .A(n2037), .ZN(n8039) );
  OAI21_X2 U12214 ( .B1(n13389), .B2(n13315), .A(n2038), .ZN(n8040) );
  OAI21_X2 U12215 ( .B1(n13484), .B2(n13315), .A(n2008), .ZN(n8041) );
  OAI21_X2 U12216 ( .B1(n13476), .B2(n13315), .A(n2009), .ZN(n8042) );
  OAI21_X2 U12217 ( .B1(n13473), .B2(n13315), .A(n2010), .ZN(n8043) );
  OAI21_X2 U12218 ( .B1(n13470), .B2(n13315), .A(n2011), .ZN(n8044) );
  OAI21_X2 U12219 ( .B1(n13467), .B2(n13315), .A(n2012), .ZN(n8045) );
  OAI21_X2 U12220 ( .B1(n13464), .B2(n13315), .A(n2013), .ZN(n8046) );
  OAI21_X2 U12221 ( .B1(n13461), .B2(n13315), .A(n2014), .ZN(n8047) );
  OAI21_X2 U12222 ( .B1(n13452), .B2(n13316), .A(n2017), .ZN(n8048) );
  OAI21_X2 U12223 ( .B1(n13419), .B2(n13317), .A(n2028), .ZN(n8049) );
  OAI21_X2 U12224 ( .B1(n13386), .B2(n13315), .A(n2039), .ZN(n8050) );
  OAI21_X2 U12225 ( .B1(n13458), .B2(n13325), .A(n1948), .ZN(n8083) );
  OAI21_X2 U12226 ( .B1(n13455), .B2(n13326), .A(n1949), .ZN(n8084) );
  OAI21_X2 U12227 ( .B1(n13449), .B2(n13326), .A(n1951), .ZN(n8085) );
  OAI21_X2 U12228 ( .B1(n13446), .B2(n13326), .A(n1952), .ZN(n8086) );
  OAI21_X2 U12229 ( .B1(n13443), .B2(n13326), .A(n1953), .ZN(n8087) );
  OAI21_X2 U12230 ( .B1(n13440), .B2(n13326), .A(n1954), .ZN(n8088) );
  OAI21_X2 U12231 ( .B1(n13437), .B2(n13326), .A(n1955), .ZN(n8089) );
  OAI21_X2 U12232 ( .B1(n13434), .B2(n13326), .A(n1956), .ZN(n8090) );
  OAI21_X2 U12233 ( .B1(n13431), .B2(n13327), .A(n1957), .ZN(n8091) );
  OAI21_X2 U12234 ( .B1(n13428), .B2(n13327), .A(n1958), .ZN(n8092) );
  OAI21_X2 U12235 ( .B1(n13425), .B2(n13326), .A(n1959), .ZN(n8093) );
  OAI21_X2 U12236 ( .B1(n13422), .B2(n13327), .A(n1960), .ZN(n8094) );
  OAI21_X2 U12237 ( .B1(n13416), .B2(n13327), .A(n1962), .ZN(n8095) );
  OAI21_X2 U12238 ( .B1(n13413), .B2(n13327), .A(n1963), .ZN(n8096) );
  OAI21_X2 U12239 ( .B1(n13410), .B2(n13327), .A(n1964), .ZN(n8097) );
  OAI21_X2 U12240 ( .B1(n13407), .B2(n13327), .A(n1965), .ZN(n8098) );
  OAI21_X2 U12241 ( .B1(n13404), .B2(n13326), .A(n1966), .ZN(n8099) );
  OAI21_X2 U12242 ( .B1(n13401), .B2(n13326), .A(n1967), .ZN(n8100) );
  OAI21_X2 U12243 ( .B1(n13398), .B2(n13326), .A(n1968), .ZN(n8101) );
  OAI21_X2 U12244 ( .B1(n13395), .B2(n13325), .A(n1969), .ZN(n8102) );
  OAI21_X2 U12245 ( .B1(n13392), .B2(n13325), .A(n1970), .ZN(n8103) );
  OAI21_X2 U12246 ( .B1(n13389), .B2(n13325), .A(n1971), .ZN(n8104) );
  OAI21_X2 U12247 ( .B1(n13484), .B2(n13325), .A(n1941), .ZN(n8105) );
  OAI21_X2 U12248 ( .B1(n13476), .B2(n13325), .A(n1942), .ZN(n8106) );
  OAI21_X2 U12249 ( .B1(n13473), .B2(n13325), .A(n1943), .ZN(n8107) );
  OAI21_X2 U12250 ( .B1(n13470), .B2(n13325), .A(n1944), .ZN(n8108) );
  OAI21_X2 U12251 ( .B1(n13467), .B2(n13325), .A(n1945), .ZN(n8109) );
  OAI21_X2 U12252 ( .B1(n13464), .B2(n13325), .A(n1946), .ZN(n8110) );
  OAI21_X2 U12253 ( .B1(n13461), .B2(n13325), .A(n1947), .ZN(n8111) );
  OAI21_X2 U12254 ( .B1(n13452), .B2(n13326), .A(n1950), .ZN(n8112) );
  OAI21_X2 U12255 ( .B1(n13419), .B2(n13327), .A(n1961), .ZN(n8113) );
  OAI21_X2 U12256 ( .B1(n13386), .B2(n13325), .A(n1972), .ZN(n8114) );
  OAI21_X2 U12257 ( .B1(n13457), .B2(n13335), .A(n1881), .ZN(n8147) );
  OAI21_X2 U12258 ( .B1(n13454), .B2(n13336), .A(n1882), .ZN(n8148) );
  OAI21_X2 U12259 ( .B1(n13448), .B2(n13336), .A(n1884), .ZN(n8149) );
  OAI21_X2 U12260 ( .B1(n13445), .B2(n13336), .A(n1885), .ZN(n8150) );
  OAI21_X2 U12261 ( .B1(n13442), .B2(n13336), .A(n1886), .ZN(n8151) );
  OAI21_X2 U12262 ( .B1(n13439), .B2(n13336), .A(n1887), .ZN(n8152) );
  OAI21_X2 U12263 ( .B1(n13436), .B2(n13336), .A(n1888), .ZN(n8153) );
  OAI21_X2 U12264 ( .B1(n13433), .B2(n13336), .A(n1889), .ZN(n8154) );
  OAI21_X2 U12265 ( .B1(n13430), .B2(n13337), .A(n1890), .ZN(n8155) );
  OAI21_X2 U12266 ( .B1(n13427), .B2(n13337), .A(n1891), .ZN(n8156) );
  OAI21_X2 U12267 ( .B1(n13424), .B2(n13336), .A(n1892), .ZN(n8157) );
  OAI21_X2 U12268 ( .B1(n13421), .B2(n13337), .A(n1893), .ZN(n8158) );
  OAI21_X2 U12269 ( .B1(n13415), .B2(n13337), .A(n1895), .ZN(n8159) );
  OAI21_X2 U12270 ( .B1(n13412), .B2(n13337), .A(n1896), .ZN(n8160) );
  OAI21_X2 U12271 ( .B1(n13409), .B2(n13337), .A(n1897), .ZN(n8161) );
  OAI21_X2 U12272 ( .B1(n13406), .B2(n13337), .A(n1898), .ZN(n8162) );
  OAI21_X2 U12273 ( .B1(n13403), .B2(n13336), .A(n1899), .ZN(n8163) );
  OAI21_X2 U12274 ( .B1(n13400), .B2(n13336), .A(n1900), .ZN(n8164) );
  OAI21_X2 U12275 ( .B1(n13397), .B2(n13336), .A(n1901), .ZN(n8165) );
  OAI21_X2 U12276 ( .B1(n13394), .B2(n13335), .A(n1902), .ZN(n8166) );
  OAI21_X2 U12277 ( .B1(n13391), .B2(n13335), .A(n1903), .ZN(n8167) );
  OAI21_X2 U12278 ( .B1(n13388), .B2(n13335), .A(n1904), .ZN(n8168) );
  OAI21_X2 U12279 ( .B1(n13483), .B2(n13335), .A(n1874), .ZN(n8169) );
  OAI21_X2 U12280 ( .B1(n13475), .B2(n13335), .A(n1875), .ZN(n8170) );
  OAI21_X2 U12281 ( .B1(n13472), .B2(n13335), .A(n1876), .ZN(n8171) );
  OAI21_X2 U12282 ( .B1(n13469), .B2(n13335), .A(n1877), .ZN(n8172) );
  OAI21_X2 U12283 ( .B1(n13466), .B2(n13335), .A(n1878), .ZN(n8173) );
  OAI21_X2 U12284 ( .B1(n13463), .B2(n13335), .A(n1879), .ZN(n8174) );
  OAI21_X2 U12285 ( .B1(n13460), .B2(n13335), .A(n1880), .ZN(n8175) );
  OAI21_X2 U12286 ( .B1(n13451), .B2(n13336), .A(n1883), .ZN(n8176) );
  OAI21_X2 U12287 ( .B1(n13418), .B2(n13337), .A(n1894), .ZN(n8177) );
  OAI21_X2 U12288 ( .B1(n13385), .B2(n13335), .A(n1905), .ZN(n8178) );
  OAI21_X2 U12289 ( .B1(n13457), .B2(n13350), .A(n1781), .ZN(n8211) );
  OAI21_X2 U12290 ( .B1(n13454), .B2(n13351), .A(n1782), .ZN(n8212) );
  OAI21_X2 U12291 ( .B1(n13448), .B2(n13351), .A(n1784), .ZN(n8213) );
  OAI21_X2 U12292 ( .B1(n13445), .B2(n13351), .A(n1785), .ZN(n8214) );
  OAI21_X2 U12293 ( .B1(n13442), .B2(n13351), .A(n1786), .ZN(n8215) );
  OAI21_X2 U12294 ( .B1(n13439), .B2(n13351), .A(n1787), .ZN(n8216) );
  OAI21_X2 U12295 ( .B1(n13436), .B2(n13351), .A(n1788), .ZN(n8217) );
  OAI21_X2 U12296 ( .B1(n13433), .B2(n13351), .A(n1789), .ZN(n8218) );
  OAI21_X2 U12297 ( .B1(n13430), .B2(n13352), .A(n1790), .ZN(n8219) );
  OAI21_X2 U12298 ( .B1(n13427), .B2(n13352), .A(n1791), .ZN(n8220) );
  OAI21_X2 U12299 ( .B1(n13424), .B2(n13351), .A(n1792), .ZN(n8221) );
  OAI21_X2 U12300 ( .B1(n13421), .B2(n13352), .A(n1793), .ZN(n8222) );
  OAI21_X2 U12301 ( .B1(n13415), .B2(n13352), .A(n1795), .ZN(n8223) );
  OAI21_X2 U12302 ( .B1(n13412), .B2(n13352), .A(n1796), .ZN(n8224) );
  OAI21_X2 U12303 ( .B1(n13409), .B2(n13352), .A(n1797), .ZN(n8225) );
  OAI21_X2 U12304 ( .B1(n13406), .B2(n13352), .A(n1798), .ZN(n8226) );
  OAI21_X2 U12305 ( .B1(n13403), .B2(n13351), .A(n1799), .ZN(n8227) );
  OAI21_X2 U12306 ( .B1(n13400), .B2(n13351), .A(n1800), .ZN(n8228) );
  OAI21_X2 U12307 ( .B1(n13397), .B2(n13351), .A(n1801), .ZN(n8229) );
  OAI21_X2 U12308 ( .B1(n13394), .B2(n13350), .A(n1802), .ZN(n8230) );
  OAI21_X2 U12309 ( .B1(n13391), .B2(n13350), .A(n1803), .ZN(n8231) );
  OAI21_X2 U12310 ( .B1(n13388), .B2(n13350), .A(n1804), .ZN(n8232) );
  OAI21_X2 U12311 ( .B1(n13483), .B2(n13350), .A(n1774), .ZN(n8233) );
  OAI21_X2 U12312 ( .B1(n13475), .B2(n13350), .A(n1775), .ZN(n8234) );
  OAI21_X2 U12313 ( .B1(n13472), .B2(n13350), .A(n1776), .ZN(n8235) );
  OAI21_X2 U12314 ( .B1(n13469), .B2(n13350), .A(n1777), .ZN(n8236) );
  OAI21_X2 U12315 ( .B1(n13466), .B2(n13350), .A(n1778), .ZN(n8237) );
  OAI21_X2 U12316 ( .B1(n13463), .B2(n13350), .A(n1779), .ZN(n8238) );
  OAI21_X2 U12317 ( .B1(n13460), .B2(n13350), .A(n1780), .ZN(n8239) );
  OAI21_X2 U12318 ( .B1(n13451), .B2(n13351), .A(n1783), .ZN(n8240) );
  OAI21_X2 U12319 ( .B1(n13418), .B2(n13352), .A(n1794), .ZN(n8241) );
  OAI21_X2 U12320 ( .B1(n13385), .B2(n13350), .A(n1805), .ZN(n8242) );
  OAI21_X2 U12321 ( .B1(n410), .B2(n13490), .A(n1480), .ZN(n6195) );
  OAI21_X2 U12322 ( .B1(n412), .B2(n13491), .A(n1481), .ZN(n6196) );
  OAI21_X2 U12323 ( .B1(n416), .B2(n13491), .A(n1483), .ZN(n6197) );
  OAI21_X2 U12324 ( .B1(n418), .B2(n13491), .A(n1484), .ZN(n6198) );
  OAI21_X2 U12325 ( .B1(n420), .B2(n13491), .A(n1485), .ZN(n6199) );
  OAI21_X2 U12326 ( .B1(n422), .B2(n13491), .A(n1486), .ZN(n6200) );
  OAI21_X2 U12327 ( .B1(n424), .B2(n13491), .A(n1487), .ZN(n6201) );
  OAI21_X2 U12328 ( .B1(n426), .B2(n13491), .A(n1488), .ZN(n6202) );
  OAI21_X2 U12329 ( .B1(n428), .B2(n13492), .A(n1489), .ZN(n6203) );
  OAI21_X2 U12330 ( .B1(n430), .B2(n13492), .A(n1490), .ZN(n6204) );
  OAI21_X2 U12331 ( .B1(n432), .B2(n13491), .A(n1491), .ZN(n6205) );
  OAI21_X2 U12332 ( .B1(n434), .B2(n13492), .A(n1492), .ZN(n6206) );
  OAI21_X2 U12333 ( .B1(n438), .B2(n13492), .A(n1494), .ZN(n6207) );
  OAI21_X2 U12334 ( .B1(n440), .B2(n13492), .A(n1495), .ZN(n6208) );
  OAI21_X2 U12335 ( .B1(n442), .B2(n13492), .A(n1496), .ZN(n6209) );
  OAI21_X2 U12336 ( .B1(n444), .B2(n13492), .A(n1497), .ZN(n6210) );
  OAI21_X2 U12337 ( .B1(n446), .B2(n13491), .A(n1498), .ZN(n6211) );
  OAI21_X2 U12338 ( .B1(n448), .B2(n13491), .A(n1499), .ZN(n6212) );
  OAI21_X2 U12339 ( .B1(n450), .B2(n13491), .A(n1500), .ZN(n6213) );
  OAI21_X2 U12340 ( .B1(n452), .B2(n13490), .A(n1501), .ZN(n6214) );
  OAI21_X2 U12341 ( .B1(n454), .B2(n13490), .A(n1502), .ZN(n6215) );
  OAI21_X2 U12342 ( .B1(n456), .B2(n13490), .A(n1503), .ZN(n6216) );
  OAI21_X2 U12343 ( .B1(n395), .B2(n13490), .A(n1471), .ZN(n6217) );
  OAI21_X2 U12344 ( .B1(n398), .B2(n13490), .A(n1474), .ZN(n6218) );
  OAI21_X2 U12345 ( .B1(n400), .B2(n13490), .A(n1475), .ZN(n6219) );
  OAI21_X2 U12346 ( .B1(n402), .B2(n13490), .A(n1476), .ZN(n6220) );
  OAI21_X2 U12347 ( .B1(n404), .B2(n13490), .A(n1477), .ZN(n6221) );
  OAI21_X2 U12348 ( .B1(n406), .B2(n13490), .A(n1478), .ZN(n6222) );
  OAI21_X2 U12349 ( .B1(n408), .B2(n13490), .A(n1479), .ZN(n6223) );
  OAI21_X2 U12350 ( .B1(n414), .B2(n13491), .A(n1482), .ZN(n6224) );
  OAI21_X2 U12351 ( .B1(n436), .B2(n13492), .A(n1493), .ZN(n6225) );
  OAI21_X2 U12352 ( .B1(n458), .B2(n13490), .A(n1504), .ZN(n6226) );
  OAI21_X2 U12353 ( .B1(n13717), .B2(n13600), .A(n742), .ZN(n6259) );
  OAI21_X2 U12354 ( .B1(n13714), .B2(n13601), .A(n743), .ZN(n6260) );
  OAI21_X2 U12355 ( .B1(n13708), .B2(n13601), .A(n745), .ZN(n6261) );
  OAI21_X2 U12356 ( .B1(n13705), .B2(n13601), .A(n746), .ZN(n6262) );
  OAI21_X2 U12357 ( .B1(n13702), .B2(n13601), .A(n747), .ZN(n6263) );
  OAI21_X2 U12358 ( .B1(n13699), .B2(n13601), .A(n748), .ZN(n6264) );
  OAI21_X2 U12359 ( .B1(n13696), .B2(n13601), .A(n749), .ZN(n6265) );
  OAI21_X2 U12360 ( .B1(n13693), .B2(n13601), .A(n750), .ZN(n6266) );
  OAI21_X2 U12361 ( .B1(n13690), .B2(n13602), .A(n751), .ZN(n6267) );
  OAI21_X2 U12362 ( .B1(n13687), .B2(n13602), .A(n752), .ZN(n6268) );
  OAI21_X2 U12363 ( .B1(n13684), .B2(n13601), .A(n753), .ZN(n6269) );
  OAI21_X2 U12364 ( .B1(n13681), .B2(n13602), .A(n754), .ZN(n6270) );
  OAI21_X2 U12365 ( .B1(n13675), .B2(n13602), .A(n756), .ZN(n6271) );
  OAI21_X2 U12366 ( .B1(n13672), .B2(n13602), .A(n757), .ZN(n6272) );
  OAI21_X2 U12367 ( .B1(n13669), .B2(n13602), .A(n758), .ZN(n6273) );
  OAI21_X2 U12368 ( .B1(n13666), .B2(n13602), .A(n759), .ZN(n6274) );
  OAI21_X2 U12369 ( .B1(n13663), .B2(n13601), .A(n760), .ZN(n6275) );
  OAI21_X2 U12370 ( .B1(n13660), .B2(n13601), .A(n761), .ZN(n6276) );
  OAI21_X2 U12371 ( .B1(n13657), .B2(n13601), .A(n762), .ZN(n6277) );
  OAI21_X2 U12372 ( .B1(n13654), .B2(n13600), .A(n763), .ZN(n6278) );
  OAI21_X2 U12373 ( .B1(n13651), .B2(n13600), .A(n764), .ZN(n6279) );
  OAI21_X2 U12374 ( .B1(n13648), .B2(n13600), .A(n765), .ZN(n6280) );
  OAI21_X2 U12375 ( .B1(n13743), .B2(n13600), .A(n735), .ZN(n6281) );
  OAI21_X2 U12376 ( .B1(n13735), .B2(n13600), .A(n736), .ZN(n6282) );
  OAI21_X2 U12377 ( .B1(n13732), .B2(n13600), .A(n737), .ZN(n6283) );
  OAI21_X2 U12378 ( .B1(n13729), .B2(n13600), .A(n738), .ZN(n6284) );
  OAI21_X2 U12379 ( .B1(n13726), .B2(n13600), .A(n739), .ZN(n6285) );
  OAI21_X2 U12380 ( .B1(n13723), .B2(n13600), .A(n740), .ZN(n6286) );
  OAI21_X2 U12381 ( .B1(n13720), .B2(n13600), .A(n741), .ZN(n6287) );
  OAI21_X2 U12382 ( .B1(n13711), .B2(n13601), .A(n744), .ZN(n6288) );
  OAI21_X2 U12383 ( .B1(n13678), .B2(n13602), .A(n755), .ZN(n6289) );
  OAI21_X2 U12384 ( .B1(n13645), .B2(n13600), .A(n766), .ZN(n6290) );
  OAI21_X2 U12385 ( .B1(n13717), .B2(n13620), .A(n606), .ZN(n6323) );
  OAI21_X2 U12386 ( .B1(n13714), .B2(n13621), .A(n607), .ZN(n6324) );
  OAI21_X2 U12387 ( .B1(n13708), .B2(n13621), .A(n609), .ZN(n6325) );
  OAI21_X2 U12388 ( .B1(n13705), .B2(n13621), .A(n610), .ZN(n6326) );
  OAI21_X2 U12389 ( .B1(n13702), .B2(n13621), .A(n611), .ZN(n6327) );
  OAI21_X2 U12390 ( .B1(n13699), .B2(n13621), .A(n612), .ZN(n6328) );
  OAI21_X2 U12391 ( .B1(n13696), .B2(n13621), .A(n613), .ZN(n6329) );
  OAI21_X2 U12392 ( .B1(n13693), .B2(n13621), .A(n614), .ZN(n6330) );
  OAI21_X2 U12393 ( .B1(n13690), .B2(n13622), .A(n615), .ZN(n6331) );
  OAI21_X2 U12394 ( .B1(n13687), .B2(n13622), .A(n616), .ZN(n6332) );
  OAI21_X2 U12395 ( .B1(n13684), .B2(n13621), .A(n617), .ZN(n6333) );
  OAI21_X2 U12396 ( .B1(n13681), .B2(n13622), .A(n618), .ZN(n6334) );
  OAI21_X2 U12397 ( .B1(n13675), .B2(n13622), .A(n620), .ZN(n6335) );
  OAI21_X2 U12398 ( .B1(n13672), .B2(n13622), .A(n621), .ZN(n6336) );
  OAI21_X2 U12399 ( .B1(n13669), .B2(n13622), .A(n622), .ZN(n6337) );
  OAI21_X2 U12400 ( .B1(n13666), .B2(n13622), .A(n623), .ZN(n6338) );
  OAI21_X2 U12401 ( .B1(n13663), .B2(n13621), .A(n624), .ZN(n6339) );
  OAI21_X2 U12402 ( .B1(n13660), .B2(n13621), .A(n625), .ZN(n6340) );
  OAI21_X2 U12403 ( .B1(n13657), .B2(n13621), .A(n626), .ZN(n6341) );
  OAI21_X2 U12404 ( .B1(n13654), .B2(n13620), .A(n627), .ZN(n6342) );
  OAI21_X2 U12405 ( .B1(n13651), .B2(n13620), .A(n628), .ZN(n6343) );
  OAI21_X2 U12406 ( .B1(n13648), .B2(n13620), .A(n629), .ZN(n6344) );
  OAI21_X2 U12407 ( .B1(n13743), .B2(n13620), .A(n599), .ZN(n6345) );
  OAI21_X2 U12408 ( .B1(n13735), .B2(n13620), .A(n600), .ZN(n6346) );
  OAI21_X2 U12409 ( .B1(n13732), .B2(n13620), .A(n601), .ZN(n6347) );
  OAI21_X2 U12410 ( .B1(n13729), .B2(n13620), .A(n602), .ZN(n6348) );
  OAI21_X2 U12411 ( .B1(n13726), .B2(n13620), .A(n603), .ZN(n6349) );
  OAI21_X2 U12412 ( .B1(n13723), .B2(n13620), .A(n604), .ZN(n6350) );
  OAI21_X2 U12413 ( .B1(n13720), .B2(n13620), .A(n605), .ZN(n6351) );
  OAI21_X2 U12414 ( .B1(n13711), .B2(n13621), .A(n608), .ZN(n6352) );
  OAI21_X2 U12415 ( .B1(n13678), .B2(n13622), .A(n619), .ZN(n6353) );
  OAI21_X2 U12416 ( .B1(n13645), .B2(n13620), .A(n630), .ZN(n6354) );
  OAI21_X2 U12417 ( .B1(n13717), .B2(n13630), .A(n539), .ZN(n6387) );
  OAI21_X2 U12418 ( .B1(n13714), .B2(n13631), .A(n540), .ZN(n6388) );
  OAI21_X2 U12419 ( .B1(n13708), .B2(n13631), .A(n542), .ZN(n6389) );
  OAI21_X2 U12420 ( .B1(n13705), .B2(n13631), .A(n543), .ZN(n6390) );
  OAI21_X2 U12421 ( .B1(n13702), .B2(n13631), .A(n544), .ZN(n6391) );
  OAI21_X2 U12422 ( .B1(n13699), .B2(n13631), .A(n545), .ZN(n6392) );
  OAI21_X2 U12423 ( .B1(n13696), .B2(n13631), .A(n546), .ZN(n6393) );
  OAI21_X2 U12424 ( .B1(n13693), .B2(n13631), .A(n547), .ZN(n6394) );
  OAI21_X2 U12425 ( .B1(n13690), .B2(n13632), .A(n548), .ZN(n6395) );
  OAI21_X2 U12426 ( .B1(n13687), .B2(n13632), .A(n549), .ZN(n6396) );
  OAI21_X2 U12427 ( .B1(n13684), .B2(n13631), .A(n550), .ZN(n6397) );
  OAI21_X2 U12428 ( .B1(n13681), .B2(n13632), .A(n551), .ZN(n6398) );
  OAI21_X2 U12429 ( .B1(n13675), .B2(n13632), .A(n553), .ZN(n6399) );
  OAI21_X2 U12430 ( .B1(n13672), .B2(n13632), .A(n554), .ZN(n6400) );
  OAI21_X2 U12431 ( .B1(n13669), .B2(n13632), .A(n555), .ZN(n6401) );
  OAI21_X2 U12432 ( .B1(n13666), .B2(n13632), .A(n556), .ZN(n6402) );
  OAI21_X2 U12433 ( .B1(n13663), .B2(n13631), .A(n557), .ZN(n6403) );
  OAI21_X2 U12434 ( .B1(n13660), .B2(n13631), .A(n558), .ZN(n6404) );
  OAI21_X2 U12435 ( .B1(n13657), .B2(n13631), .A(n559), .ZN(n6405) );
  OAI21_X2 U12436 ( .B1(n13654), .B2(n13630), .A(n560), .ZN(n6406) );
  OAI21_X2 U12437 ( .B1(n13651), .B2(n13630), .A(n561), .ZN(n6407) );
  OAI21_X2 U12438 ( .B1(n13648), .B2(n13630), .A(n562), .ZN(n6408) );
  OAI21_X2 U12439 ( .B1(n13743), .B2(n13630), .A(n532), .ZN(n6409) );
  OAI21_X2 U12440 ( .B1(n13735), .B2(n13630), .A(n533), .ZN(n6410) );
  OAI21_X2 U12441 ( .B1(n13732), .B2(n13630), .A(n534), .ZN(n6411) );
  OAI21_X2 U12442 ( .B1(n13729), .B2(n13630), .A(n535), .ZN(n6412) );
  OAI21_X2 U12443 ( .B1(n13726), .B2(n13630), .A(n536), .ZN(n6413) );
  OAI21_X2 U12444 ( .B1(n13723), .B2(n13630), .A(n537), .ZN(n6414) );
  OAI21_X2 U12445 ( .B1(n13720), .B2(n13630), .A(n538), .ZN(n6415) );
  OAI21_X2 U12446 ( .B1(n13711), .B2(n13631), .A(n541), .ZN(n6416) );
  OAI21_X2 U12447 ( .B1(n13678), .B2(n13632), .A(n552), .ZN(n6417) );
  OAI21_X2 U12448 ( .B1(n13645), .B2(n13630), .A(n563), .ZN(n6418) );
  OAI21_X2 U12449 ( .B1(n13717), .B2(n13640), .A(n470), .ZN(n6451) );
  OAI21_X2 U12450 ( .B1(n13714), .B2(n13641), .A(n471), .ZN(n6452) );
  OAI21_X2 U12451 ( .B1(n13708), .B2(n13641), .A(n473), .ZN(n6453) );
  OAI21_X2 U12452 ( .B1(n13705), .B2(n13641), .A(n474), .ZN(n6454) );
  OAI21_X2 U12453 ( .B1(n13702), .B2(n13641), .A(n475), .ZN(n6455) );
  OAI21_X2 U12454 ( .B1(n13699), .B2(n13641), .A(n476), .ZN(n6456) );
  OAI21_X2 U12455 ( .B1(n13696), .B2(n13641), .A(n477), .ZN(n6457) );
  OAI21_X2 U12456 ( .B1(n13693), .B2(n13641), .A(n478), .ZN(n6458) );
  OAI21_X2 U12457 ( .B1(n13690), .B2(n13642), .A(n479), .ZN(n6459) );
  OAI21_X2 U12458 ( .B1(n13687), .B2(n13642), .A(n480), .ZN(n6460) );
  OAI21_X2 U12459 ( .B1(n13684), .B2(n13641), .A(n481), .ZN(n6461) );
  OAI21_X2 U12460 ( .B1(n13681), .B2(n13642), .A(n482), .ZN(n6462) );
  OAI21_X2 U12461 ( .B1(n13675), .B2(n13642), .A(n484), .ZN(n6463) );
  OAI21_X2 U12462 ( .B1(n13672), .B2(n13642), .A(n485), .ZN(n6464) );
  OAI21_X2 U12463 ( .B1(n13669), .B2(n13642), .A(n486), .ZN(n6465) );
  OAI21_X2 U12464 ( .B1(n13666), .B2(n13642), .A(n487), .ZN(n6466) );
  OAI21_X2 U12465 ( .B1(n13663), .B2(n13641), .A(n488), .ZN(n6467) );
  OAI21_X2 U12466 ( .B1(n13660), .B2(n13641), .A(n489), .ZN(n6468) );
  OAI21_X2 U12467 ( .B1(n13657), .B2(n13641), .A(n490), .ZN(n6469) );
  OAI21_X2 U12468 ( .B1(n13654), .B2(n13640), .A(n491), .ZN(n6470) );
  OAI21_X2 U12469 ( .B1(n13651), .B2(n13640), .A(n492), .ZN(n6471) );
  OAI21_X2 U12470 ( .B1(n13648), .B2(n13640), .A(n493), .ZN(n6472) );
  OAI21_X2 U12471 ( .B1(n13743), .B2(n13640), .A(n463), .ZN(n6473) );
  OAI21_X2 U12472 ( .B1(n13735), .B2(n13640), .A(n464), .ZN(n6474) );
  OAI21_X2 U12473 ( .B1(n13732), .B2(n13640), .A(n465), .ZN(n6475) );
  OAI21_X2 U12474 ( .B1(n13729), .B2(n13640), .A(n466), .ZN(n6476) );
  OAI21_X2 U12475 ( .B1(n13726), .B2(n13640), .A(n467), .ZN(n6477) );
  OAI21_X2 U12476 ( .B1(n13723), .B2(n13640), .A(n468), .ZN(n6478) );
  OAI21_X2 U12477 ( .B1(n13720), .B2(n13640), .A(n469), .ZN(n6479) );
  OAI21_X2 U12478 ( .B1(n13711), .B2(n13641), .A(n472), .ZN(n6480) );
  OAI21_X2 U12479 ( .B1(n13678), .B2(n13642), .A(n483), .ZN(n6481) );
  OAI21_X2 U12480 ( .B1(n13645), .B2(n13640), .A(n494), .ZN(n6482) );
  OAI21_X2 U12481 ( .B1(n410), .B2(n13495), .A(n1445), .ZN(n6515) );
  OAI21_X2 U12482 ( .B1(n412), .B2(n13496), .A(n1446), .ZN(n6516) );
  OAI21_X2 U12483 ( .B1(n416), .B2(n13496), .A(n1448), .ZN(n6517) );
  OAI21_X2 U12484 ( .B1(n418), .B2(n13496), .A(n1449), .ZN(n6518) );
  OAI21_X2 U12485 ( .B1(n420), .B2(n13496), .A(n1450), .ZN(n6519) );
  OAI21_X2 U12486 ( .B1(n422), .B2(n13496), .A(n1451), .ZN(n6520) );
  OAI21_X2 U12487 ( .B1(n424), .B2(n13496), .A(n1452), .ZN(n6521) );
  OAI21_X2 U12488 ( .B1(n426), .B2(n13496), .A(n1453), .ZN(n6522) );
  OAI21_X2 U12489 ( .B1(n428), .B2(n13497), .A(n1454), .ZN(n6523) );
  OAI21_X2 U12490 ( .B1(n430), .B2(n13497), .A(n1455), .ZN(n6524) );
  OAI21_X2 U12491 ( .B1(n432), .B2(n13496), .A(n1456), .ZN(n6525) );
  OAI21_X2 U12492 ( .B1(n434), .B2(n13497), .A(n1457), .ZN(n6526) );
  OAI21_X2 U12493 ( .B1(n438), .B2(n13497), .A(n1459), .ZN(n6527) );
  OAI21_X2 U12494 ( .B1(n440), .B2(n13497), .A(n1460), .ZN(n6528) );
  OAI21_X2 U12495 ( .B1(n442), .B2(n13497), .A(n1461), .ZN(n6529) );
  OAI21_X2 U12496 ( .B1(n444), .B2(n13497), .A(n1462), .ZN(n6530) );
  OAI21_X2 U12497 ( .B1(n446), .B2(n13496), .A(n1463), .ZN(n6531) );
  OAI21_X2 U12498 ( .B1(n448), .B2(n13496), .A(n1464), .ZN(n6532) );
  OAI21_X2 U12499 ( .B1(n450), .B2(n13496), .A(n1465), .ZN(n6533) );
  OAI21_X2 U12500 ( .B1(n452), .B2(n13495), .A(n1466), .ZN(n6534) );
  OAI21_X2 U12501 ( .B1(n454), .B2(n13495), .A(n1467), .ZN(n6535) );
  OAI21_X2 U12502 ( .B1(n456), .B2(n13495), .A(n1468), .ZN(n6536) );
  OAI21_X2 U12503 ( .B1(n395), .B2(n13495), .A(n1438), .ZN(n6537) );
  OAI21_X2 U12504 ( .B1(n398), .B2(n13495), .A(n1439), .ZN(n6538) );
  OAI21_X2 U12505 ( .B1(n400), .B2(n13495), .A(n1440), .ZN(n6539) );
  OAI21_X2 U12506 ( .B1(n402), .B2(n13495), .A(n1441), .ZN(n6540) );
  OAI21_X2 U12507 ( .B1(n404), .B2(n13495), .A(n1442), .ZN(n6541) );
  OAI21_X2 U12508 ( .B1(n406), .B2(n13495), .A(n1443), .ZN(n6542) );
  OAI21_X2 U12509 ( .B1(n408), .B2(n13495), .A(n1444), .ZN(n6543) );
  OAI21_X2 U12510 ( .B1(n414), .B2(n13496), .A(n1447), .ZN(n6544) );
  OAI21_X2 U12511 ( .B1(n436), .B2(n13497), .A(n1458), .ZN(n6545) );
  OAI21_X2 U12512 ( .B1(n458), .B2(n13495), .A(n1469), .ZN(n6546) );
  OAI21_X2 U12513 ( .B1(n410), .B2(n13505), .A(n1379), .ZN(n6579) );
  OAI21_X2 U12514 ( .B1(n412), .B2(n13506), .A(n1380), .ZN(n6580) );
  OAI21_X2 U12515 ( .B1(n416), .B2(n13506), .A(n1382), .ZN(n6581) );
  OAI21_X2 U12516 ( .B1(n418), .B2(n13506), .A(n1383), .ZN(n6582) );
  OAI21_X2 U12517 ( .B1(n420), .B2(n13506), .A(n1384), .ZN(n6583) );
  OAI21_X2 U12518 ( .B1(n422), .B2(n13506), .A(n1385), .ZN(n6584) );
  OAI21_X2 U12519 ( .B1(n424), .B2(n13506), .A(n1386), .ZN(n6585) );
  OAI21_X2 U12520 ( .B1(n426), .B2(n13506), .A(n1387), .ZN(n6586) );
  OAI21_X2 U12521 ( .B1(n428), .B2(n13507), .A(n1388), .ZN(n6587) );
  OAI21_X2 U12522 ( .B1(n430), .B2(n13507), .A(n1389), .ZN(n6588) );
  OAI21_X2 U12523 ( .B1(n432), .B2(n13506), .A(n1390), .ZN(n6589) );
  OAI21_X2 U12524 ( .B1(n434), .B2(n13507), .A(n1391), .ZN(n6590) );
  OAI21_X2 U12525 ( .B1(n438), .B2(n13507), .A(n1393), .ZN(n6591) );
  OAI21_X2 U12526 ( .B1(n440), .B2(n13507), .A(n1394), .ZN(n6592) );
  OAI21_X2 U12527 ( .B1(n442), .B2(n13507), .A(n1395), .ZN(n6593) );
  OAI21_X2 U12528 ( .B1(n444), .B2(n13507), .A(n1396), .ZN(n6594) );
  OAI21_X2 U12529 ( .B1(n446), .B2(n13506), .A(n1397), .ZN(n6595) );
  OAI21_X2 U12530 ( .B1(n448), .B2(n13506), .A(n1398), .ZN(n6596) );
  OAI21_X2 U12531 ( .B1(n450), .B2(n13506), .A(n1399), .ZN(n6597) );
  OAI21_X2 U12532 ( .B1(n452), .B2(n13505), .A(n1400), .ZN(n6598) );
  OAI21_X2 U12533 ( .B1(n454), .B2(n13505), .A(n1401), .ZN(n6599) );
  OAI21_X2 U12534 ( .B1(n456), .B2(n13505), .A(n1402), .ZN(n6600) );
  OAI21_X2 U12535 ( .B1(n395), .B2(n13505), .A(n1372), .ZN(n6601) );
  OAI21_X2 U12536 ( .B1(n398), .B2(n13505), .A(n1373), .ZN(n6602) );
  OAI21_X2 U12537 ( .B1(n400), .B2(n13505), .A(n1374), .ZN(n6603) );
  OAI21_X2 U12538 ( .B1(n402), .B2(n13505), .A(n1375), .ZN(n6604) );
  OAI21_X2 U12539 ( .B1(n404), .B2(n13505), .A(n1376), .ZN(n6605) );
  OAI21_X2 U12540 ( .B1(n406), .B2(n13505), .A(n1377), .ZN(n6606) );
  OAI21_X2 U12541 ( .B1(n408), .B2(n13505), .A(n1378), .ZN(n6607) );
  OAI21_X2 U12542 ( .B1(n414), .B2(n13506), .A(n1381), .ZN(n6608) );
  OAI21_X2 U12543 ( .B1(n436), .B2(n13507), .A(n1392), .ZN(n6609) );
  OAI21_X2 U12544 ( .B1(n458), .B2(n13505), .A(n1403), .ZN(n6610) );
  OAI21_X2 U12545 ( .B1(n410), .B2(n13515), .A(n1312), .ZN(n6643) );
  OAI21_X2 U12546 ( .B1(n412), .B2(n13516), .A(n1313), .ZN(n6644) );
  OAI21_X2 U12547 ( .B1(n416), .B2(n13516), .A(n1315), .ZN(n6645) );
  OAI21_X2 U12548 ( .B1(n418), .B2(n13516), .A(n1316), .ZN(n6646) );
  OAI21_X2 U12549 ( .B1(n420), .B2(n13516), .A(n1317), .ZN(n6647) );
  OAI21_X2 U12550 ( .B1(n422), .B2(n13516), .A(n1318), .ZN(n6648) );
  OAI21_X2 U12551 ( .B1(n424), .B2(n13516), .A(n1319), .ZN(n6649) );
  OAI21_X2 U12552 ( .B1(n426), .B2(n13516), .A(n1320), .ZN(n6650) );
  OAI21_X2 U12553 ( .B1(n428), .B2(n13517), .A(n1321), .ZN(n6651) );
  OAI21_X2 U12554 ( .B1(n430), .B2(n13517), .A(n1322), .ZN(n6652) );
  OAI21_X2 U12555 ( .B1(n432), .B2(n13516), .A(n1323), .ZN(n6653) );
  OAI21_X2 U12556 ( .B1(n434), .B2(n13517), .A(n1324), .ZN(n6654) );
  OAI21_X2 U12557 ( .B1(n438), .B2(n13517), .A(n1326), .ZN(n6655) );
  OAI21_X2 U12558 ( .B1(n440), .B2(n13517), .A(n1327), .ZN(n6656) );
  OAI21_X2 U12559 ( .B1(n442), .B2(n13517), .A(n1328), .ZN(n6657) );
  OAI21_X2 U12560 ( .B1(n444), .B2(n13517), .A(n1329), .ZN(n6658) );
  OAI21_X2 U12561 ( .B1(n446), .B2(n13516), .A(n1330), .ZN(n6659) );
  OAI21_X2 U12562 ( .B1(n448), .B2(n13516), .A(n1331), .ZN(n6660) );
  OAI21_X2 U12563 ( .B1(n450), .B2(n13516), .A(n1332), .ZN(n6661) );
  OAI21_X2 U12564 ( .B1(n452), .B2(n13515), .A(n1333), .ZN(n6662) );
  OAI21_X2 U12565 ( .B1(n454), .B2(n13515), .A(n1334), .ZN(n6663) );
  OAI21_X2 U12566 ( .B1(n456), .B2(n13515), .A(n1335), .ZN(n6664) );
  OAI21_X2 U12567 ( .B1(n395), .B2(n13515), .A(n1305), .ZN(n6665) );
  OAI21_X2 U12568 ( .B1(n398), .B2(n13515), .A(n1306), .ZN(n6666) );
  OAI21_X2 U12569 ( .B1(n400), .B2(n13515), .A(n1307), .ZN(n6667) );
  OAI21_X2 U12570 ( .B1(n402), .B2(n13515), .A(n1308), .ZN(n6668) );
  OAI21_X2 U12571 ( .B1(n404), .B2(n13515), .A(n1309), .ZN(n6669) );
  OAI21_X2 U12572 ( .B1(n406), .B2(n13515), .A(n1310), .ZN(n6670) );
  OAI21_X2 U12573 ( .B1(n408), .B2(n13515), .A(n1311), .ZN(n6671) );
  OAI21_X2 U12574 ( .B1(n414), .B2(n13516), .A(n1314), .ZN(n6672) );
  OAI21_X2 U12575 ( .B1(n436), .B2(n13517), .A(n1325), .ZN(n6673) );
  OAI21_X2 U12576 ( .B1(n458), .B2(n13515), .A(n1336), .ZN(n6674) );
  OAI21_X2 U12577 ( .B1(n410), .B2(n13525), .A(n1244), .ZN(n6707) );
  OAI21_X2 U12578 ( .B1(n412), .B2(n13526), .A(n1245), .ZN(n6708) );
  OAI21_X2 U12579 ( .B1(n416), .B2(n13526), .A(n1247), .ZN(n6709) );
  OAI21_X2 U12580 ( .B1(n418), .B2(n13526), .A(n1248), .ZN(n6710) );
  OAI21_X2 U12581 ( .B1(n420), .B2(n13526), .A(n1249), .ZN(n6711) );
  OAI21_X2 U12582 ( .B1(n422), .B2(n13526), .A(n1250), .ZN(n6712) );
  OAI21_X2 U12583 ( .B1(n424), .B2(n13526), .A(n1251), .ZN(n6713) );
  OAI21_X2 U12584 ( .B1(n426), .B2(n13526), .A(n1252), .ZN(n6714) );
  OAI21_X2 U12585 ( .B1(n428), .B2(n13527), .A(n1253), .ZN(n6715) );
  OAI21_X2 U12586 ( .B1(n430), .B2(n13527), .A(n1254), .ZN(n6716) );
  OAI21_X2 U12587 ( .B1(n432), .B2(n13526), .A(n1255), .ZN(n6717) );
  OAI21_X2 U12588 ( .B1(n434), .B2(n13527), .A(n1256), .ZN(n6718) );
  OAI21_X2 U12589 ( .B1(n438), .B2(n13527), .A(n1258), .ZN(n6719) );
  OAI21_X2 U12590 ( .B1(n440), .B2(n13527), .A(n1259), .ZN(n6720) );
  OAI21_X2 U12591 ( .B1(n442), .B2(n13527), .A(n1260), .ZN(n6721) );
  OAI21_X2 U12592 ( .B1(n444), .B2(n13527), .A(n1261), .ZN(n6722) );
  OAI21_X2 U12593 ( .B1(n446), .B2(n13526), .A(n1262), .ZN(n6723) );
  OAI21_X2 U12594 ( .B1(n448), .B2(n13526), .A(n1263), .ZN(n6724) );
  OAI21_X2 U12595 ( .B1(n450), .B2(n13526), .A(n1264), .ZN(n6725) );
  OAI21_X2 U12596 ( .B1(n452), .B2(n13525), .A(n1265), .ZN(n6726) );
  OAI21_X2 U12597 ( .B1(n454), .B2(n13525), .A(n1266), .ZN(n6727) );
  OAI21_X2 U12598 ( .B1(n456), .B2(n13525), .A(n1267), .ZN(n6728) );
  OAI21_X2 U12599 ( .B1(n395), .B2(n13525), .A(n1237), .ZN(n6729) );
  OAI21_X2 U12600 ( .B1(n398), .B2(n13525), .A(n1238), .ZN(n6730) );
  OAI21_X2 U12601 ( .B1(n400), .B2(n13525), .A(n1239), .ZN(n6731) );
  OAI21_X2 U12602 ( .B1(n402), .B2(n13525), .A(n1240), .ZN(n6732) );
  OAI21_X2 U12603 ( .B1(n404), .B2(n13525), .A(n1241), .ZN(n6733) );
  OAI21_X2 U12604 ( .B1(n406), .B2(n13525), .A(n1242), .ZN(n6734) );
  OAI21_X2 U12605 ( .B1(n408), .B2(n13525), .A(n1243), .ZN(n6735) );
  OAI21_X2 U12606 ( .B1(n414), .B2(n13526), .A(n1246), .ZN(n6736) );
  OAI21_X2 U12607 ( .B1(n436), .B2(n13527), .A(n1257), .ZN(n6737) );
  OAI21_X2 U12608 ( .B1(n458), .B2(n13525), .A(n1268), .ZN(n6738) );
  OAI21_X2 U12609 ( .B1(n13718), .B2(n13535), .A(n1178), .ZN(n6771) );
  OAI21_X2 U12610 ( .B1(n13715), .B2(n13536), .A(n1179), .ZN(n6772) );
  OAI21_X2 U12611 ( .B1(n13709), .B2(n13536), .A(n1181), .ZN(n6773) );
  OAI21_X2 U12612 ( .B1(n13706), .B2(n13536), .A(n1182), .ZN(n6774) );
  OAI21_X2 U12613 ( .B1(n13703), .B2(n13536), .A(n1183), .ZN(n6775) );
  OAI21_X2 U12614 ( .B1(n13700), .B2(n13536), .A(n1184), .ZN(n6776) );
  OAI21_X2 U12615 ( .B1(n13697), .B2(n13536), .A(n1185), .ZN(n6777) );
  OAI21_X2 U12616 ( .B1(n13694), .B2(n13536), .A(n1186), .ZN(n6778) );
  OAI21_X2 U12617 ( .B1(n13691), .B2(n13537), .A(n1187), .ZN(n6779) );
  OAI21_X2 U12618 ( .B1(n13688), .B2(n13537), .A(n1188), .ZN(n6780) );
  OAI21_X2 U12619 ( .B1(n13685), .B2(n13536), .A(n1189), .ZN(n6781) );
  OAI21_X2 U12620 ( .B1(n13682), .B2(n13537), .A(n1190), .ZN(n6782) );
  OAI21_X2 U12621 ( .B1(n13676), .B2(n13537), .A(n1192), .ZN(n6783) );
  OAI21_X2 U12622 ( .B1(n13673), .B2(n13537), .A(n1193), .ZN(n6784) );
  OAI21_X2 U12623 ( .B1(n13670), .B2(n13537), .A(n1194), .ZN(n6785) );
  OAI21_X2 U12624 ( .B1(n13667), .B2(n13537), .A(n1195), .ZN(n6786) );
  OAI21_X2 U12625 ( .B1(n13664), .B2(n13536), .A(n1196), .ZN(n6787) );
  OAI21_X2 U12626 ( .B1(n13661), .B2(n13536), .A(n1197), .ZN(n6788) );
  OAI21_X2 U12627 ( .B1(n13658), .B2(n13536), .A(n1198), .ZN(n6789) );
  OAI21_X2 U12628 ( .B1(n13655), .B2(n13535), .A(n1199), .ZN(n6790) );
  OAI21_X2 U12629 ( .B1(n13652), .B2(n13535), .A(n1200), .ZN(n6791) );
  OAI21_X2 U12630 ( .B1(n13649), .B2(n13535), .A(n1201), .ZN(n6792) );
  OAI21_X2 U12631 ( .B1(n13744), .B2(n13535), .A(n1171), .ZN(n6793) );
  OAI21_X2 U12632 ( .B1(n13736), .B2(n13535), .A(n1172), .ZN(n6794) );
  OAI21_X2 U12633 ( .B1(n13733), .B2(n13535), .A(n1173), .ZN(n6795) );
  OAI21_X2 U12634 ( .B1(n13730), .B2(n13535), .A(n1174), .ZN(n6796) );
  OAI21_X2 U12635 ( .B1(n13727), .B2(n13535), .A(n1175), .ZN(n6797) );
  OAI21_X2 U12636 ( .B1(n13724), .B2(n13535), .A(n1176), .ZN(n6798) );
  OAI21_X2 U12637 ( .B1(n13721), .B2(n13535), .A(n1177), .ZN(n6799) );
  OAI21_X2 U12638 ( .B1(n13712), .B2(n13536), .A(n1180), .ZN(n6800) );
  OAI21_X2 U12639 ( .B1(n13679), .B2(n13537), .A(n1191), .ZN(n6801) );
  OAI21_X2 U12640 ( .B1(n13646), .B2(n13535), .A(n1202), .ZN(n6802) );
  OAI21_X2 U12641 ( .B1(n13718), .B2(n13550), .A(n1078), .ZN(n6835) );
  OAI21_X2 U12642 ( .B1(n13715), .B2(n13551), .A(n1079), .ZN(n6836) );
  OAI21_X2 U12643 ( .B1(n13709), .B2(n13551), .A(n1081), .ZN(n6837) );
  OAI21_X2 U12644 ( .B1(n13706), .B2(n13551), .A(n1082), .ZN(n6838) );
  OAI21_X2 U12645 ( .B1(n13703), .B2(n13551), .A(n1083), .ZN(n6839) );
  OAI21_X2 U12646 ( .B1(n13700), .B2(n13551), .A(n1084), .ZN(n6840) );
  OAI21_X2 U12647 ( .B1(n13697), .B2(n13551), .A(n1085), .ZN(n6841) );
  OAI21_X2 U12648 ( .B1(n13694), .B2(n13551), .A(n1086), .ZN(n6842) );
  OAI21_X2 U12649 ( .B1(n13691), .B2(n13552), .A(n1087), .ZN(n6843) );
  OAI21_X2 U12650 ( .B1(n13688), .B2(n13552), .A(n1088), .ZN(n6844) );
  OAI21_X2 U12651 ( .B1(n13685), .B2(n13551), .A(n1089), .ZN(n6845) );
  OAI21_X2 U12652 ( .B1(n13682), .B2(n13552), .A(n1090), .ZN(n6846) );
  OAI21_X2 U12653 ( .B1(n13676), .B2(n13552), .A(n1092), .ZN(n6847) );
  OAI21_X2 U12654 ( .B1(n13673), .B2(n13552), .A(n1093), .ZN(n6848) );
  OAI21_X2 U12655 ( .B1(n13670), .B2(n13552), .A(n1094), .ZN(n6849) );
  OAI21_X2 U12656 ( .B1(n13667), .B2(n13552), .A(n1095), .ZN(n6850) );
  OAI21_X2 U12657 ( .B1(n13664), .B2(n13551), .A(n1096), .ZN(n6851) );
  OAI21_X2 U12658 ( .B1(n13661), .B2(n13551), .A(n1097), .ZN(n6852) );
  OAI21_X2 U12659 ( .B1(n13658), .B2(n13551), .A(n1098), .ZN(n6853) );
  OAI21_X2 U12660 ( .B1(n13655), .B2(n13550), .A(n1099), .ZN(n6854) );
  OAI21_X2 U12661 ( .B1(n13652), .B2(n13550), .A(n1100), .ZN(n6855) );
  OAI21_X2 U12662 ( .B1(n13649), .B2(n13550), .A(n1101), .ZN(n6856) );
  OAI21_X2 U12663 ( .B1(n13744), .B2(n13550), .A(n1071), .ZN(n6857) );
  OAI21_X2 U12664 ( .B1(n13736), .B2(n13550), .A(n1072), .ZN(n6858) );
  OAI21_X2 U12665 ( .B1(n13733), .B2(n13550), .A(n1073), .ZN(n6859) );
  OAI21_X2 U12666 ( .B1(n13730), .B2(n13550), .A(n1074), .ZN(n6860) );
  OAI21_X2 U12667 ( .B1(n13727), .B2(n13550), .A(n1075), .ZN(n6861) );
  OAI21_X2 U12668 ( .B1(n13724), .B2(n13550), .A(n1076), .ZN(n6862) );
  OAI21_X2 U12669 ( .B1(n13721), .B2(n13550), .A(n1077), .ZN(n6863) );
  OAI21_X2 U12670 ( .B1(n13712), .B2(n13551), .A(n1080), .ZN(n6864) );
  OAI21_X2 U12671 ( .B1(n13679), .B2(n13552), .A(n1091), .ZN(n6865) );
  OAI21_X2 U12672 ( .B1(n13646), .B2(n13550), .A(n1102), .ZN(n6866) );
  OAI21_X2 U12673 ( .B1(n13718), .B2(n13560), .A(n1012), .ZN(n6899) );
  OAI21_X2 U12674 ( .B1(n13715), .B2(n13561), .A(n1013), .ZN(n6900) );
  OAI21_X2 U12675 ( .B1(n13709), .B2(n13561), .A(n1015), .ZN(n6901) );
  OAI21_X2 U12676 ( .B1(n13706), .B2(n13561), .A(n1016), .ZN(n6902) );
  OAI21_X2 U12677 ( .B1(n13703), .B2(n13561), .A(n1017), .ZN(n6903) );
  OAI21_X2 U12678 ( .B1(n13700), .B2(n13561), .A(n1018), .ZN(n6904) );
  OAI21_X2 U12679 ( .B1(n13697), .B2(n13561), .A(n1019), .ZN(n6905) );
  OAI21_X2 U12680 ( .B1(n13694), .B2(n13561), .A(n1020), .ZN(n6906) );
  OAI21_X2 U12681 ( .B1(n13691), .B2(n13562), .A(n1021), .ZN(n6907) );
  OAI21_X2 U12682 ( .B1(n13688), .B2(n13562), .A(n1022), .ZN(n6908) );
  OAI21_X2 U12683 ( .B1(n13685), .B2(n13561), .A(n1023), .ZN(n6909) );
  OAI21_X2 U12684 ( .B1(n13682), .B2(n13562), .A(n1024), .ZN(n6910) );
  OAI21_X2 U12685 ( .B1(n13676), .B2(n13562), .A(n1026), .ZN(n6911) );
  OAI21_X2 U12686 ( .B1(n13673), .B2(n13562), .A(n1027), .ZN(n6912) );
  OAI21_X2 U12687 ( .B1(n13670), .B2(n13562), .A(n1028), .ZN(n6913) );
  OAI21_X2 U12688 ( .B1(n13667), .B2(n13562), .A(n1029), .ZN(n6914) );
  OAI21_X2 U12689 ( .B1(n13664), .B2(n13561), .A(n1030), .ZN(n6915) );
  OAI21_X2 U12690 ( .B1(n13661), .B2(n13561), .A(n1031), .ZN(n6916) );
  OAI21_X2 U12691 ( .B1(n13658), .B2(n13561), .A(n1032), .ZN(n6917) );
  OAI21_X2 U12692 ( .B1(n13655), .B2(n13560), .A(n1033), .ZN(n6918) );
  OAI21_X2 U12693 ( .B1(n13652), .B2(n13560), .A(n1034), .ZN(n6919) );
  OAI21_X2 U12694 ( .B1(n13649), .B2(n13560), .A(n1035), .ZN(n6920) );
  OAI21_X2 U12695 ( .B1(n13744), .B2(n13560), .A(n1005), .ZN(n6921) );
  OAI21_X2 U12696 ( .B1(n13736), .B2(n13560), .A(n1006), .ZN(n6922) );
  OAI21_X2 U12697 ( .B1(n13733), .B2(n13560), .A(n1007), .ZN(n6923) );
  OAI21_X2 U12698 ( .B1(n13730), .B2(n13560), .A(n1008), .ZN(n6924) );
  OAI21_X2 U12699 ( .B1(n13727), .B2(n13560), .A(n1009), .ZN(n6925) );
  OAI21_X2 U12700 ( .B1(n13724), .B2(n13560), .A(n1010), .ZN(n6926) );
  OAI21_X2 U12701 ( .B1(n13721), .B2(n13560), .A(n1011), .ZN(n6927) );
  OAI21_X2 U12702 ( .B1(n13712), .B2(n13561), .A(n1014), .ZN(n6928) );
  OAI21_X2 U12703 ( .B1(n13679), .B2(n13562), .A(n1025), .ZN(n6929) );
  OAI21_X2 U12704 ( .B1(n13646), .B2(n13560), .A(n1036), .ZN(n6930) );
  OAI21_X2 U12705 ( .B1(n13718), .B2(n13570), .A(n945), .ZN(n6963) );
  OAI21_X2 U12706 ( .B1(n13715), .B2(n13571), .A(n946), .ZN(n6964) );
  OAI21_X2 U12707 ( .B1(n13709), .B2(n13571), .A(n948), .ZN(n6965) );
  OAI21_X2 U12708 ( .B1(n13706), .B2(n13571), .A(n949), .ZN(n6966) );
  OAI21_X2 U12709 ( .B1(n13703), .B2(n13571), .A(n950), .ZN(n6967) );
  OAI21_X2 U12710 ( .B1(n13700), .B2(n13571), .A(n951), .ZN(n6968) );
  OAI21_X2 U12711 ( .B1(n13697), .B2(n13571), .A(n952), .ZN(n6969) );
  OAI21_X2 U12712 ( .B1(n13694), .B2(n13571), .A(n953), .ZN(n6970) );
  OAI21_X2 U12713 ( .B1(n13691), .B2(n13572), .A(n954), .ZN(n6971) );
  OAI21_X2 U12714 ( .B1(n13688), .B2(n13572), .A(n955), .ZN(n6972) );
  OAI21_X2 U12715 ( .B1(n13685), .B2(n13571), .A(n956), .ZN(n6973) );
  OAI21_X2 U12716 ( .B1(n13682), .B2(n13572), .A(n957), .ZN(n6974) );
  OAI21_X2 U12717 ( .B1(n13676), .B2(n13572), .A(n959), .ZN(n6975) );
  OAI21_X2 U12718 ( .B1(n13673), .B2(n13572), .A(n960), .ZN(n6976) );
  OAI21_X2 U12719 ( .B1(n13670), .B2(n13572), .A(n961), .ZN(n6977) );
  OAI21_X2 U12720 ( .B1(n13667), .B2(n13572), .A(n962), .ZN(n6978) );
  OAI21_X2 U12721 ( .B1(n13664), .B2(n13571), .A(n963), .ZN(n6979) );
  OAI21_X2 U12722 ( .B1(n13661), .B2(n13571), .A(n964), .ZN(n6980) );
  OAI21_X2 U12723 ( .B1(n13658), .B2(n13571), .A(n965), .ZN(n6981) );
  OAI21_X2 U12724 ( .B1(n13655), .B2(n13570), .A(n966), .ZN(n6982) );
  OAI21_X2 U12725 ( .B1(n13652), .B2(n13570), .A(n967), .ZN(n6983) );
  OAI21_X2 U12726 ( .B1(n13649), .B2(n13570), .A(n968), .ZN(n6984) );
  OAI21_X2 U12727 ( .B1(n13744), .B2(n13570), .A(n938), .ZN(n6985) );
  OAI21_X2 U12728 ( .B1(n13736), .B2(n13570), .A(n939), .ZN(n6986) );
  OAI21_X2 U12729 ( .B1(n13733), .B2(n13570), .A(n940), .ZN(n6987) );
  OAI21_X2 U12730 ( .B1(n13730), .B2(n13570), .A(n941), .ZN(n6988) );
  OAI21_X2 U12731 ( .B1(n13727), .B2(n13570), .A(n942), .ZN(n6989) );
  OAI21_X2 U12732 ( .B1(n13724), .B2(n13570), .A(n943), .ZN(n6990) );
  OAI21_X2 U12733 ( .B1(n13721), .B2(n13570), .A(n944), .ZN(n6991) );
  OAI21_X2 U12734 ( .B1(n13712), .B2(n13571), .A(n947), .ZN(n6992) );
  OAI21_X2 U12735 ( .B1(n13679), .B2(n13572), .A(n958), .ZN(n6993) );
  OAI21_X2 U12736 ( .B1(n13646), .B2(n13570), .A(n969), .ZN(n6994) );
  OAI21_X2 U12737 ( .B1(n13718), .B2(n13580), .A(n879), .ZN(n7027) );
  OAI21_X2 U12738 ( .B1(n13715), .B2(n13581), .A(n880), .ZN(n7028) );
  OAI21_X2 U12739 ( .B1(n13709), .B2(n13581), .A(n882), .ZN(n7029) );
  OAI21_X2 U12740 ( .B1(n13706), .B2(n13581), .A(n883), .ZN(n7030) );
  OAI21_X2 U12741 ( .B1(n13703), .B2(n13581), .A(n884), .ZN(n7031) );
  OAI21_X2 U12742 ( .B1(n13700), .B2(n13581), .A(n885), .ZN(n7032) );
  OAI21_X2 U12743 ( .B1(n13697), .B2(n13581), .A(n886), .ZN(n7033) );
  OAI21_X2 U12744 ( .B1(n13694), .B2(n13581), .A(n887), .ZN(n7034) );
  OAI21_X2 U12745 ( .B1(n13691), .B2(n13582), .A(n888), .ZN(n7035) );
  OAI21_X2 U12746 ( .B1(n13688), .B2(n13582), .A(n889), .ZN(n7036) );
  OAI21_X2 U12747 ( .B1(n13685), .B2(n13581), .A(n890), .ZN(n7037) );
  OAI21_X2 U12748 ( .B1(n13682), .B2(n13582), .A(n891), .ZN(n7038) );
  OAI21_X2 U12749 ( .B1(n13676), .B2(n13582), .A(n893), .ZN(n7039) );
  OAI21_X2 U12750 ( .B1(n13673), .B2(n13582), .A(n894), .ZN(n7040) );
  OAI21_X2 U12751 ( .B1(n13670), .B2(n13582), .A(n895), .ZN(n7041) );
  OAI21_X2 U12752 ( .B1(n13667), .B2(n13582), .A(n896), .ZN(n7042) );
  OAI21_X2 U12753 ( .B1(n13664), .B2(n13581), .A(n897), .ZN(n7043) );
  OAI21_X2 U12754 ( .B1(n13661), .B2(n13581), .A(n898), .ZN(n7044) );
  OAI21_X2 U12755 ( .B1(n13658), .B2(n13581), .A(n899), .ZN(n7045) );
  OAI21_X2 U12756 ( .B1(n13655), .B2(n13580), .A(n900), .ZN(n7046) );
  OAI21_X2 U12757 ( .B1(n13652), .B2(n13580), .A(n901), .ZN(n7047) );
  OAI21_X2 U12758 ( .B1(n13649), .B2(n13580), .A(n902), .ZN(n7048) );
  OAI21_X2 U12759 ( .B1(n13744), .B2(n13580), .A(n872), .ZN(n7049) );
  OAI21_X2 U12760 ( .B1(n13736), .B2(n13580), .A(n873), .ZN(n7050) );
  OAI21_X2 U12761 ( .B1(n13733), .B2(n13580), .A(n874), .ZN(n7051) );
  OAI21_X2 U12762 ( .B1(n13730), .B2(n13580), .A(n875), .ZN(n7052) );
  OAI21_X2 U12763 ( .B1(n13727), .B2(n13580), .A(n876), .ZN(n7053) );
  OAI21_X2 U12764 ( .B1(n13724), .B2(n13580), .A(n877), .ZN(n7054) );
  OAI21_X2 U12765 ( .B1(n13721), .B2(n13580), .A(n878), .ZN(n7055) );
  OAI21_X2 U12766 ( .B1(n13712), .B2(n13581), .A(n881), .ZN(n7056) );
  OAI21_X2 U12767 ( .B1(n13679), .B2(n13582), .A(n892), .ZN(n7057) );
  OAI21_X2 U12768 ( .B1(n13646), .B2(n13580), .A(n903), .ZN(n7058) );
  OAI21_X2 U12769 ( .B1(n13717), .B2(n13590), .A(n809), .ZN(n7091) );
  OAI21_X2 U12770 ( .B1(n13714), .B2(n13591), .A(n810), .ZN(n7092) );
  OAI21_X2 U12771 ( .B1(n13708), .B2(n13591), .A(n812), .ZN(n7093) );
  OAI21_X2 U12772 ( .B1(n13705), .B2(n13591), .A(n813), .ZN(n7094) );
  OAI21_X2 U12773 ( .B1(n13702), .B2(n13591), .A(n814), .ZN(n7095) );
  OAI21_X2 U12774 ( .B1(n13699), .B2(n13591), .A(n815), .ZN(n7096) );
  OAI21_X2 U12775 ( .B1(n13696), .B2(n13591), .A(n816), .ZN(n7097) );
  OAI21_X2 U12776 ( .B1(n13693), .B2(n13591), .A(n817), .ZN(n7098) );
  OAI21_X2 U12777 ( .B1(n13690), .B2(n13592), .A(n818), .ZN(n7099) );
  OAI21_X2 U12778 ( .B1(n13687), .B2(n13592), .A(n819), .ZN(n7100) );
  OAI21_X2 U12779 ( .B1(n13684), .B2(n13591), .A(n820), .ZN(n7101) );
  OAI21_X2 U12780 ( .B1(n13681), .B2(n13592), .A(n821), .ZN(n7102) );
  OAI21_X2 U12781 ( .B1(n13675), .B2(n13592), .A(n823), .ZN(n7103) );
  OAI21_X2 U12782 ( .B1(n13672), .B2(n13592), .A(n824), .ZN(n7104) );
  OAI21_X2 U12783 ( .B1(n13669), .B2(n13592), .A(n825), .ZN(n7105) );
  OAI21_X2 U12784 ( .B1(n13666), .B2(n13592), .A(n826), .ZN(n7106) );
  OAI21_X2 U12785 ( .B1(n13663), .B2(n13591), .A(n827), .ZN(n7107) );
  OAI21_X2 U12786 ( .B1(n13660), .B2(n13591), .A(n828), .ZN(n7108) );
  OAI21_X2 U12787 ( .B1(n13657), .B2(n13591), .A(n829), .ZN(n7109) );
  OAI21_X2 U12788 ( .B1(n13654), .B2(n13590), .A(n830), .ZN(n7110) );
  OAI21_X2 U12789 ( .B1(n13651), .B2(n13590), .A(n831), .ZN(n7111) );
  OAI21_X2 U12790 ( .B1(n13648), .B2(n13590), .A(n832), .ZN(n7112) );
  OAI21_X2 U12791 ( .B1(n13743), .B2(n13590), .A(n802), .ZN(n7113) );
  OAI21_X2 U12792 ( .B1(n13735), .B2(n13590), .A(n803), .ZN(n7114) );
  OAI21_X2 U12793 ( .B1(n13732), .B2(n13590), .A(n804), .ZN(n7115) );
  OAI21_X2 U12794 ( .B1(n13729), .B2(n13590), .A(n805), .ZN(n7116) );
  OAI21_X2 U12795 ( .B1(n13726), .B2(n13590), .A(n806), .ZN(n7117) );
  OAI21_X2 U12796 ( .B1(n13723), .B2(n13590), .A(n807), .ZN(n7118) );
  OAI21_X2 U12797 ( .B1(n13720), .B2(n13590), .A(n808), .ZN(n7119) );
  OAI21_X2 U12798 ( .B1(n13711), .B2(n13591), .A(n811), .ZN(n7120) );
  OAI21_X2 U12799 ( .B1(n13678), .B2(n13592), .A(n822), .ZN(n7121) );
  OAI21_X2 U12800 ( .B1(n13645), .B2(n13590), .A(n833), .ZN(n7122) );
  OAI21_X2 U12801 ( .B1(n13717), .B2(n13605), .A(n708), .ZN(n7155) );
  OAI21_X2 U12802 ( .B1(n13714), .B2(n13606), .A(n709), .ZN(n7156) );
  OAI21_X2 U12803 ( .B1(n13708), .B2(n13606), .A(n711), .ZN(n7157) );
  OAI21_X2 U12804 ( .B1(n13705), .B2(n13606), .A(n712), .ZN(n7158) );
  OAI21_X2 U12805 ( .B1(n13702), .B2(n13606), .A(n713), .ZN(n7159) );
  OAI21_X2 U12806 ( .B1(n13699), .B2(n13606), .A(n714), .ZN(n7160) );
  OAI21_X2 U12807 ( .B1(n13696), .B2(n13606), .A(n715), .ZN(n7161) );
  OAI21_X2 U12808 ( .B1(n13693), .B2(n13606), .A(n716), .ZN(n7162) );
  OAI21_X2 U12809 ( .B1(n13690), .B2(n13607), .A(n717), .ZN(n7163) );
  OAI21_X2 U12810 ( .B1(n13687), .B2(n13607), .A(n718), .ZN(n7164) );
  OAI21_X2 U12811 ( .B1(n13684), .B2(n13606), .A(n719), .ZN(n7165) );
  OAI21_X2 U12812 ( .B1(n13681), .B2(n13607), .A(n720), .ZN(n7166) );
  OAI21_X2 U12813 ( .B1(n13675), .B2(n13607), .A(n722), .ZN(n7167) );
  OAI21_X2 U12814 ( .B1(n13672), .B2(n13607), .A(n723), .ZN(n7168) );
  OAI21_X2 U12815 ( .B1(n13669), .B2(n13607), .A(n724), .ZN(n7169) );
  OAI21_X2 U12816 ( .B1(n13666), .B2(n13607), .A(n725), .ZN(n7170) );
  OAI21_X2 U12817 ( .B1(n13663), .B2(n13606), .A(n726), .ZN(n7171) );
  OAI21_X2 U12818 ( .B1(n13660), .B2(n13606), .A(n727), .ZN(n7172) );
  OAI21_X2 U12819 ( .B1(n13657), .B2(n13606), .A(n728), .ZN(n7173) );
  OAI21_X2 U12820 ( .B1(n13654), .B2(n13605), .A(n729), .ZN(n7174) );
  OAI21_X2 U12821 ( .B1(n13651), .B2(n13605), .A(n730), .ZN(n7175) );
  OAI21_X2 U12822 ( .B1(n13648), .B2(n13605), .A(n731), .ZN(n7176) );
  OAI21_X2 U12823 ( .B1(n13743), .B2(n13605), .A(n701), .ZN(n7177) );
  OAI21_X2 U12824 ( .B1(n13735), .B2(n13605), .A(n702), .ZN(n7178) );
  OAI21_X2 U12825 ( .B1(n13732), .B2(n13605), .A(n703), .ZN(n7179) );
  OAI21_X2 U12826 ( .B1(n13729), .B2(n13605), .A(n704), .ZN(n7180) );
  OAI21_X2 U12827 ( .B1(n13726), .B2(n13605), .A(n705), .ZN(n7181) );
  OAI21_X2 U12828 ( .B1(n13723), .B2(n13605), .A(n706), .ZN(n7182) );
  OAI21_X2 U12829 ( .B1(n13720), .B2(n13605), .A(n707), .ZN(n7183) );
  OAI21_X2 U12830 ( .B1(n13711), .B2(n13606), .A(n710), .ZN(n7184) );
  OAI21_X2 U12831 ( .B1(n13678), .B2(n13607), .A(n721), .ZN(n7185) );
  OAI21_X2 U12832 ( .B1(n13645), .B2(n13605), .A(n732), .ZN(n7186) );
  OAI21_X2 U12833 ( .B1(n1521), .B2(n13230), .A(n2592), .ZN(n7219) );
  OAI21_X2 U12834 ( .B1(n1523), .B2(n13231), .A(n2594), .ZN(n7220) );
  OAI21_X2 U12835 ( .B1(n1527), .B2(n13231), .A(n2598), .ZN(n7221) );
  OAI21_X2 U12836 ( .B1(n1529), .B2(n13231), .A(n2600), .ZN(n7222) );
  OAI21_X2 U12837 ( .B1(n1531), .B2(n13231), .A(n2602), .ZN(n7223) );
  OAI21_X2 U12838 ( .B1(n1533), .B2(n13231), .A(n2604), .ZN(n7224) );
  OAI21_X2 U12839 ( .B1(n1535), .B2(n13231), .A(n2606), .ZN(n7225) );
  OAI21_X2 U12840 ( .B1(n1537), .B2(n13231), .A(n2608), .ZN(n7226) );
  OAI21_X2 U12841 ( .B1(n1539), .B2(n13232), .A(n2610), .ZN(n7227) );
  OAI21_X2 U12842 ( .B1(n1541), .B2(n13232), .A(n2612), .ZN(n7228) );
  OAI21_X2 U12843 ( .B1(n1543), .B2(n13231), .A(n2614), .ZN(n7229) );
  OAI21_X2 U12844 ( .B1(n1545), .B2(n13232), .A(n2616), .ZN(n7230) );
  OAI21_X2 U12845 ( .B1(n1549), .B2(n13232), .A(n2620), .ZN(n7231) );
  OAI21_X2 U12846 ( .B1(n1551), .B2(n13232), .A(n2622), .ZN(n7232) );
  OAI21_X2 U12847 ( .B1(n1553), .B2(n13232), .A(n2624), .ZN(n7233) );
  OAI21_X2 U12848 ( .B1(n1555), .B2(n13232), .A(n2626), .ZN(n7234) );
  OAI21_X2 U12849 ( .B1(n1557), .B2(n13231), .A(n2628), .ZN(n7235) );
  OAI21_X2 U12850 ( .B1(n1559), .B2(n13231), .A(n2630), .ZN(n7236) );
  OAI21_X2 U12851 ( .B1(n1561), .B2(n13231), .A(n2632), .ZN(n7237) );
  OAI21_X2 U12852 ( .B1(n1563), .B2(n13230), .A(n2634), .ZN(n7238) );
  OAI21_X2 U12853 ( .B1(n1565), .B2(n13230), .A(n2636), .ZN(n7239) );
  OAI21_X2 U12854 ( .B1(n1567), .B2(n13230), .A(n2638), .ZN(n7240) );
  OAI21_X2 U12855 ( .B1(n1506), .B2(n13230), .A(n2576), .ZN(n7241) );
  OAI21_X2 U12856 ( .B1(n1509), .B2(n13230), .A(n2580), .ZN(n7242) );
  OAI21_X2 U12857 ( .B1(n1511), .B2(n13230), .A(n2582), .ZN(n7243) );
  OAI21_X2 U12858 ( .B1(n1513), .B2(n13230), .A(n2584), .ZN(n7244) );
  OAI21_X2 U12859 ( .B1(n1515), .B2(n13230), .A(n2586), .ZN(n7245) );
  OAI21_X2 U12860 ( .B1(n1517), .B2(n13230), .A(n2588), .ZN(n7246) );
  OAI21_X2 U12861 ( .B1(n1519), .B2(n13230), .A(n2590), .ZN(n7247) );
  OAI21_X2 U12862 ( .B1(n1525), .B2(n13231), .A(n2596), .ZN(n7248) );
  OAI21_X2 U12863 ( .B1(n1547), .B2(n13232), .A(n2618), .ZN(n7249) );
  OAI21_X2 U12864 ( .B1(n1569), .B2(n13230), .A(n2640), .ZN(n7250) );
  OAI21_X2 U12865 ( .B1(n13457), .B2(n13340), .A(n1848), .ZN(n7283) );
  OAI21_X2 U12866 ( .B1(n13454), .B2(n13341), .A(n1849), .ZN(n7284) );
  OAI21_X2 U12867 ( .B1(n13448), .B2(n13341), .A(n1851), .ZN(n7285) );
  OAI21_X2 U12868 ( .B1(n13445), .B2(n13341), .A(n1852), .ZN(n7286) );
  OAI21_X2 U12869 ( .B1(n13442), .B2(n13341), .A(n1853), .ZN(n7287) );
  OAI21_X2 U12870 ( .B1(n13439), .B2(n13341), .A(n1854), .ZN(n7288) );
  OAI21_X2 U12871 ( .B1(n13436), .B2(n13341), .A(n1855), .ZN(n7289) );
  OAI21_X2 U12872 ( .B1(n13433), .B2(n13341), .A(n1856), .ZN(n7290) );
  OAI21_X2 U12873 ( .B1(n13430), .B2(n13342), .A(n1857), .ZN(n7291) );
  OAI21_X2 U12874 ( .B1(n13427), .B2(n13342), .A(n1858), .ZN(n7292) );
  OAI21_X2 U12875 ( .B1(n13424), .B2(n13341), .A(n1859), .ZN(n7293) );
  OAI21_X2 U12876 ( .B1(n13421), .B2(n13342), .A(n1860), .ZN(n7294) );
  OAI21_X2 U12877 ( .B1(n13415), .B2(n13342), .A(n1862), .ZN(n7295) );
  OAI21_X2 U12878 ( .B1(n13412), .B2(n13342), .A(n1863), .ZN(n7296) );
  OAI21_X2 U12879 ( .B1(n13409), .B2(n13342), .A(n1864), .ZN(n7297) );
  OAI21_X2 U12880 ( .B1(n13406), .B2(n13342), .A(n1865), .ZN(n7298) );
  OAI21_X2 U12881 ( .B1(n13403), .B2(n13341), .A(n1866), .ZN(n7299) );
  OAI21_X2 U12882 ( .B1(n13400), .B2(n13341), .A(n1867), .ZN(n7300) );
  OAI21_X2 U12883 ( .B1(n13397), .B2(n13341), .A(n1868), .ZN(n7301) );
  OAI21_X2 U12884 ( .B1(n13394), .B2(n13340), .A(n1869), .ZN(n7302) );
  OAI21_X2 U12885 ( .B1(n13391), .B2(n13340), .A(n1870), .ZN(n7303) );
  OAI21_X2 U12886 ( .B1(n13388), .B2(n13340), .A(n1871), .ZN(n7304) );
  OAI21_X2 U12887 ( .B1(n13483), .B2(n13340), .A(n1841), .ZN(n7305) );
  OAI21_X2 U12888 ( .B1(n13475), .B2(n13340), .A(n1842), .ZN(n7306) );
  OAI21_X2 U12889 ( .B1(n13472), .B2(n13340), .A(n1843), .ZN(n7307) );
  OAI21_X2 U12890 ( .B1(n13469), .B2(n13340), .A(n1844), .ZN(n7308) );
  OAI21_X2 U12891 ( .B1(n13466), .B2(n13340), .A(n1845), .ZN(n7309) );
  OAI21_X2 U12892 ( .B1(n13463), .B2(n13340), .A(n1846), .ZN(n7310) );
  OAI21_X2 U12893 ( .B1(n13460), .B2(n13340), .A(n1847), .ZN(n7311) );
  OAI21_X2 U12894 ( .B1(n13451), .B2(n13341), .A(n1850), .ZN(n7312) );
  OAI21_X2 U12895 ( .B1(n13418), .B2(n13342), .A(n1861), .ZN(n7313) );
  OAI21_X2 U12896 ( .B1(n13385), .B2(n13340), .A(n1872), .ZN(n7314) );
  OAI21_X2 U12897 ( .B1(n13457), .B2(n13360), .A(n1713), .ZN(n7347) );
  OAI21_X2 U12898 ( .B1(n13454), .B2(n13361), .A(n1714), .ZN(n7348) );
  OAI21_X2 U12899 ( .B1(n13448), .B2(n13361), .A(n1716), .ZN(n7349) );
  OAI21_X2 U12900 ( .B1(n13445), .B2(n13361), .A(n1717), .ZN(n7350) );
  OAI21_X2 U12901 ( .B1(n13442), .B2(n13361), .A(n1718), .ZN(n7351) );
  OAI21_X2 U12902 ( .B1(n13439), .B2(n13361), .A(n1719), .ZN(n7352) );
  OAI21_X2 U12903 ( .B1(n13436), .B2(n13361), .A(n1720), .ZN(n7353) );
  OAI21_X2 U12904 ( .B1(n13433), .B2(n13361), .A(n1721), .ZN(n7354) );
  OAI21_X2 U12905 ( .B1(n13430), .B2(n13362), .A(n1722), .ZN(n7355) );
  OAI21_X2 U12906 ( .B1(n13427), .B2(n13362), .A(n1723), .ZN(n7356) );
  OAI21_X2 U12907 ( .B1(n13424), .B2(n13361), .A(n1724), .ZN(n7357) );
  OAI21_X2 U12908 ( .B1(n13421), .B2(n13362), .A(n1725), .ZN(n7358) );
  OAI21_X2 U12909 ( .B1(n13415), .B2(n13362), .A(n1727), .ZN(n7359) );
  OAI21_X2 U12910 ( .B1(n13412), .B2(n13362), .A(n1728), .ZN(n7360) );
  OAI21_X2 U12911 ( .B1(n13409), .B2(n13362), .A(n1729), .ZN(n7361) );
  OAI21_X2 U12912 ( .B1(n13406), .B2(n13362), .A(n1730), .ZN(n7362) );
  OAI21_X2 U12913 ( .B1(n13403), .B2(n13361), .A(n1731), .ZN(n7363) );
  OAI21_X2 U12914 ( .B1(n13400), .B2(n13361), .A(n1732), .ZN(n7364) );
  OAI21_X2 U12915 ( .B1(n13397), .B2(n13361), .A(n1733), .ZN(n7365) );
  OAI21_X2 U12916 ( .B1(n13394), .B2(n13360), .A(n1734), .ZN(n7366) );
  OAI21_X2 U12917 ( .B1(n13391), .B2(n13360), .A(n1735), .ZN(n7367) );
  OAI21_X2 U12918 ( .B1(n13388), .B2(n13360), .A(n1736), .ZN(n7368) );
  OAI21_X2 U12919 ( .B1(n13483), .B2(n13360), .A(n1706), .ZN(n7369) );
  OAI21_X2 U12920 ( .B1(n13475), .B2(n13360), .A(n1707), .ZN(n7370) );
  OAI21_X2 U12921 ( .B1(n13472), .B2(n13360), .A(n1708), .ZN(n7371) );
  OAI21_X2 U12922 ( .B1(n13469), .B2(n13360), .A(n1709), .ZN(n7372) );
  OAI21_X2 U12923 ( .B1(n13466), .B2(n13360), .A(n1710), .ZN(n7373) );
  OAI21_X2 U12924 ( .B1(n13463), .B2(n13360), .A(n1711), .ZN(n7374) );
  OAI21_X2 U12925 ( .B1(n13460), .B2(n13360), .A(n1712), .ZN(n7375) );
  OAI21_X2 U12926 ( .B1(n13451), .B2(n13361), .A(n1715), .ZN(n7376) );
  OAI21_X2 U12927 ( .B1(n13418), .B2(n13362), .A(n1726), .ZN(n7377) );
  OAI21_X2 U12928 ( .B1(n13385), .B2(n13360), .A(n1737), .ZN(n7378) );
  OAI21_X2 U12929 ( .B1(n13457), .B2(n13370), .A(n1647), .ZN(n7411) );
  OAI21_X2 U12930 ( .B1(n13454), .B2(n13371), .A(n1648), .ZN(n7412) );
  OAI21_X2 U12931 ( .B1(n13448), .B2(n13371), .A(n1650), .ZN(n7413) );
  OAI21_X2 U12932 ( .B1(n13445), .B2(n13371), .A(n1651), .ZN(n7414) );
  OAI21_X2 U12933 ( .B1(n13442), .B2(n13371), .A(n1652), .ZN(n7415) );
  OAI21_X2 U12934 ( .B1(n13439), .B2(n13371), .A(n1653), .ZN(n7416) );
  OAI21_X2 U12935 ( .B1(n13436), .B2(n13371), .A(n1654), .ZN(n7417) );
  OAI21_X2 U12936 ( .B1(n13433), .B2(n13371), .A(n1655), .ZN(n7418) );
  OAI21_X2 U12937 ( .B1(n13430), .B2(n13372), .A(n1656), .ZN(n7419) );
  OAI21_X2 U12938 ( .B1(n13427), .B2(n13372), .A(n1657), .ZN(n7420) );
  OAI21_X2 U12939 ( .B1(n13424), .B2(n13371), .A(n1658), .ZN(n7421) );
  OAI21_X2 U12940 ( .B1(n13421), .B2(n13372), .A(n1659), .ZN(n7422) );
  OAI21_X2 U12941 ( .B1(n13415), .B2(n13372), .A(n1661), .ZN(n7423) );
  OAI21_X2 U12942 ( .B1(n13412), .B2(n13372), .A(n1662), .ZN(n7424) );
  OAI21_X2 U12943 ( .B1(n13409), .B2(n13372), .A(n1663), .ZN(n7425) );
  OAI21_X2 U12944 ( .B1(n13406), .B2(n13372), .A(n1664), .ZN(n7426) );
  OAI21_X2 U12945 ( .B1(n13403), .B2(n13371), .A(n1665), .ZN(n7427) );
  OAI21_X2 U12946 ( .B1(n13400), .B2(n13371), .A(n1666), .ZN(n7428) );
  OAI21_X2 U12947 ( .B1(n13397), .B2(n13371), .A(n1667), .ZN(n7429) );
  OAI21_X2 U12948 ( .B1(n13394), .B2(n13370), .A(n1668), .ZN(n7430) );
  OAI21_X2 U12949 ( .B1(n13391), .B2(n13370), .A(n1669), .ZN(n7431) );
  OAI21_X2 U12950 ( .B1(n13388), .B2(n13370), .A(n1670), .ZN(n7432) );
  OAI21_X2 U12951 ( .B1(n13483), .B2(n13370), .A(n1640), .ZN(n7433) );
  OAI21_X2 U12952 ( .B1(n13475), .B2(n13370), .A(n1641), .ZN(n7434) );
  OAI21_X2 U12953 ( .B1(n13472), .B2(n13370), .A(n1642), .ZN(n7435) );
  OAI21_X2 U12954 ( .B1(n13469), .B2(n13370), .A(n1643), .ZN(n7436) );
  OAI21_X2 U12955 ( .B1(n13466), .B2(n13370), .A(n1644), .ZN(n7437) );
  OAI21_X2 U12956 ( .B1(n13463), .B2(n13370), .A(n1645), .ZN(n7438) );
  OAI21_X2 U12957 ( .B1(n13460), .B2(n13370), .A(n1646), .ZN(n7439) );
  OAI21_X2 U12958 ( .B1(n13451), .B2(n13371), .A(n1649), .ZN(n7440) );
  OAI21_X2 U12959 ( .B1(n13418), .B2(n13372), .A(n1660), .ZN(n7441) );
  OAI21_X2 U12960 ( .B1(n13385), .B2(n13370), .A(n1671), .ZN(n7442) );
  OAI21_X2 U12961 ( .B1(n13457), .B2(n13380), .A(n1580), .ZN(n7475) );
  OAI21_X2 U12962 ( .B1(n13454), .B2(n13381), .A(n1581), .ZN(n7476) );
  OAI21_X2 U12963 ( .B1(n13448), .B2(n13381), .A(n1583), .ZN(n7477) );
  OAI21_X2 U12964 ( .B1(n13445), .B2(n13381), .A(n1584), .ZN(n7478) );
  OAI21_X2 U12965 ( .B1(n13442), .B2(n13381), .A(n1585), .ZN(n7479) );
  OAI21_X2 U12966 ( .B1(n13439), .B2(n13381), .A(n1586), .ZN(n7480) );
  OAI21_X2 U12967 ( .B1(n13436), .B2(n13381), .A(n1587), .ZN(n7481) );
  OAI21_X2 U12968 ( .B1(n13433), .B2(n13381), .A(n1588), .ZN(n7482) );
  OAI21_X2 U12969 ( .B1(n13430), .B2(n13382), .A(n1589), .ZN(n7483) );
  OAI21_X2 U12970 ( .B1(n13427), .B2(n13382), .A(n1590), .ZN(n7484) );
  OAI21_X2 U12971 ( .B1(n13424), .B2(n13381), .A(n1591), .ZN(n7485) );
  OAI21_X2 U12972 ( .B1(n13421), .B2(n13382), .A(n1592), .ZN(n7486) );
  OAI21_X2 U12973 ( .B1(n13415), .B2(n13382), .A(n1594), .ZN(n7487) );
  OAI21_X2 U12974 ( .B1(n13412), .B2(n13382), .A(n1595), .ZN(n7488) );
  OAI21_X2 U12975 ( .B1(n13409), .B2(n13382), .A(n1596), .ZN(n7489) );
  OAI21_X2 U12976 ( .B1(n13406), .B2(n13382), .A(n1597), .ZN(n7490) );
  OAI21_X2 U12977 ( .B1(n13403), .B2(n13381), .A(n1598), .ZN(n7491) );
  OAI21_X2 U12978 ( .B1(n13400), .B2(n13381), .A(n1599), .ZN(n7492) );
  OAI21_X2 U12979 ( .B1(n13397), .B2(n13381), .A(n1600), .ZN(n7493) );
  OAI21_X2 U12980 ( .B1(n13394), .B2(n13380), .A(n1601), .ZN(n7494) );
  OAI21_X2 U12981 ( .B1(n13391), .B2(n13380), .A(n1602), .ZN(n7495) );
  OAI21_X2 U12982 ( .B1(n13388), .B2(n13380), .A(n1603), .ZN(n7496) );
  OAI21_X2 U12983 ( .B1(n13483), .B2(n13380), .A(n1573), .ZN(n7497) );
  OAI21_X2 U12984 ( .B1(n13475), .B2(n13380), .A(n1574), .ZN(n7498) );
  OAI21_X2 U12985 ( .B1(n13472), .B2(n13380), .A(n1575), .ZN(n7499) );
  OAI21_X2 U12986 ( .B1(n13469), .B2(n13380), .A(n1576), .ZN(n7500) );
  OAI21_X2 U12987 ( .B1(n13466), .B2(n13380), .A(n1577), .ZN(n7501) );
  OAI21_X2 U12988 ( .B1(n13463), .B2(n13380), .A(n1578), .ZN(n7502) );
  OAI21_X2 U12989 ( .B1(n13460), .B2(n13380), .A(n1579), .ZN(n7503) );
  OAI21_X2 U12990 ( .B1(n13451), .B2(n13381), .A(n1582), .ZN(n7504) );
  OAI21_X2 U12991 ( .B1(n13418), .B2(n13382), .A(n1593), .ZN(n7505) );
  OAI21_X2 U12992 ( .B1(n13385), .B2(n13380), .A(n1604), .ZN(n7506) );
  OAI21_X2 U12993 ( .B1(n1521), .B2(n13235), .A(n2550), .ZN(n7539) );
  OAI21_X2 U12994 ( .B1(n1523), .B2(n13236), .A(n2551), .ZN(n7540) );
  OAI21_X2 U12995 ( .B1(n1527), .B2(n13236), .A(n2553), .ZN(n7541) );
  OAI21_X2 U12996 ( .B1(n1529), .B2(n13236), .A(n2554), .ZN(n7542) );
  OAI21_X2 U12997 ( .B1(n1531), .B2(n13236), .A(n2555), .ZN(n7543) );
  OAI21_X2 U12998 ( .B1(n1533), .B2(n13236), .A(n2556), .ZN(n7544) );
  OAI21_X2 U12999 ( .B1(n1535), .B2(n13236), .A(n2557), .ZN(n7545) );
  OAI21_X2 U13000 ( .B1(n1537), .B2(n13236), .A(n2558), .ZN(n7546) );
  OAI21_X2 U13001 ( .B1(n1539), .B2(n13237), .A(n2559), .ZN(n7547) );
  OAI21_X2 U13002 ( .B1(n1541), .B2(n13237), .A(n2560), .ZN(n7548) );
  OAI21_X2 U13003 ( .B1(n1543), .B2(n13236), .A(n2561), .ZN(n7549) );
  OAI21_X2 U13004 ( .B1(n1545), .B2(n13237), .A(n2562), .ZN(n7550) );
  OAI21_X2 U13005 ( .B1(n1549), .B2(n13237), .A(n2564), .ZN(n7551) );
  OAI21_X2 U13006 ( .B1(n1551), .B2(n13237), .A(n2565), .ZN(n7552) );
  OAI21_X2 U13007 ( .B1(n1553), .B2(n13237), .A(n2566), .ZN(n7553) );
  OAI21_X2 U13008 ( .B1(n1555), .B2(n13237), .A(n2567), .ZN(n7554) );
  OAI21_X2 U13009 ( .B1(n1557), .B2(n13236), .A(n2568), .ZN(n7555) );
  OAI21_X2 U13010 ( .B1(n1559), .B2(n13236), .A(n2569), .ZN(n7556) );
  OAI21_X2 U13011 ( .B1(n1561), .B2(n13236), .A(n2570), .ZN(n7557) );
  OAI21_X2 U13012 ( .B1(n1563), .B2(n13235), .A(n2571), .ZN(n7558) );
  OAI21_X2 U13013 ( .B1(n1565), .B2(n13235), .A(n2572), .ZN(n7559) );
  OAI21_X2 U13014 ( .B1(n1567), .B2(n13235), .A(n2573), .ZN(n7560) );
  OAI21_X2 U13015 ( .B1(n1506), .B2(n13235), .A(n2543), .ZN(n7561) );
  OAI21_X2 U13016 ( .B1(n1509), .B2(n13235), .A(n2544), .ZN(n7562) );
  OAI21_X2 U13017 ( .B1(n1511), .B2(n13235), .A(n2545), .ZN(n7563) );
  OAI21_X2 U13018 ( .B1(n1513), .B2(n13235), .A(n2546), .ZN(n7564) );
  OAI21_X2 U13019 ( .B1(n1515), .B2(n13235), .A(n2547), .ZN(n7565) );
  OAI21_X2 U13020 ( .B1(n1517), .B2(n13235), .A(n2548), .ZN(n7566) );
  OAI21_X2 U13021 ( .B1(n1519), .B2(n13235), .A(n2549), .ZN(n7567) );
  OAI21_X2 U13022 ( .B1(n1525), .B2(n13236), .A(n2552), .ZN(n7568) );
  OAI21_X2 U13023 ( .B1(n1547), .B2(n13237), .A(n2563), .ZN(n7569) );
  OAI21_X2 U13024 ( .B1(n1569), .B2(n13235), .A(n2574), .ZN(n7570) );
  OAI21_X2 U13025 ( .B1(n1521), .B2(n13245), .A(n2483), .ZN(n7603) );
  OAI21_X2 U13026 ( .B1(n1523), .B2(n13246), .A(n2484), .ZN(n7604) );
  OAI21_X2 U13027 ( .B1(n1527), .B2(n13246), .A(n2486), .ZN(n7605) );
  OAI21_X2 U13028 ( .B1(n1529), .B2(n13246), .A(n2487), .ZN(n7606) );
  OAI21_X2 U13029 ( .B1(n1531), .B2(n13246), .A(n2488), .ZN(n7607) );
  OAI21_X2 U13030 ( .B1(n1533), .B2(n13246), .A(n2489), .ZN(n7608) );
  OAI21_X2 U13031 ( .B1(n1535), .B2(n13246), .A(n2490), .ZN(n7609) );
  OAI21_X2 U13032 ( .B1(n1537), .B2(n13246), .A(n2491), .ZN(n7610) );
  OAI21_X2 U13033 ( .B1(n1539), .B2(n13247), .A(n2492), .ZN(n7611) );
  OAI21_X2 U13034 ( .B1(n1541), .B2(n13247), .A(n2493), .ZN(n7612) );
  OAI21_X2 U13035 ( .B1(n1543), .B2(n13246), .A(n2494), .ZN(n7613) );
  OAI21_X2 U13036 ( .B1(n1545), .B2(n13247), .A(n2495), .ZN(n7614) );
  OAI21_X2 U13037 ( .B1(n1549), .B2(n13247), .A(n2497), .ZN(n7615) );
  OAI21_X2 U13038 ( .B1(n1551), .B2(n13247), .A(n2498), .ZN(n7616) );
  OAI21_X2 U13039 ( .B1(n1553), .B2(n13247), .A(n2499), .ZN(n7617) );
  OAI21_X2 U13040 ( .B1(n1555), .B2(n13247), .A(n2500), .ZN(n7618) );
  OAI21_X2 U13041 ( .B1(n1557), .B2(n13246), .A(n2501), .ZN(n7619) );
  OAI21_X2 U13042 ( .B1(n1559), .B2(n13246), .A(n2502), .ZN(n7620) );
  OAI21_X2 U13043 ( .B1(n1561), .B2(n13246), .A(n2503), .ZN(n7621) );
  OAI21_X2 U13044 ( .B1(n1563), .B2(n13245), .A(n2504), .ZN(n7622) );
  OAI21_X2 U13045 ( .B1(n1565), .B2(n13245), .A(n2505), .ZN(n7623) );
  OAI21_X2 U13046 ( .B1(n1567), .B2(n13245), .A(n2506), .ZN(n7624) );
  OAI21_X2 U13047 ( .B1(n1506), .B2(n13245), .A(n2476), .ZN(n7625) );
  OAI21_X2 U13048 ( .B1(n1509), .B2(n13245), .A(n2477), .ZN(n7626) );
  OAI21_X2 U13049 ( .B1(n1511), .B2(n13245), .A(n2478), .ZN(n7627) );
  OAI21_X2 U13050 ( .B1(n1513), .B2(n13245), .A(n2479), .ZN(n7628) );
  OAI21_X2 U13051 ( .B1(n1515), .B2(n13245), .A(n2480), .ZN(n7629) );
  OAI21_X2 U13052 ( .B1(n1517), .B2(n13245), .A(n2481), .ZN(n7630) );
  OAI21_X2 U13053 ( .B1(n1519), .B2(n13245), .A(n2482), .ZN(n7631) );
  OAI21_X2 U13054 ( .B1(n1525), .B2(n13246), .A(n2485), .ZN(n7632) );
  OAI21_X2 U13055 ( .B1(n1547), .B2(n13247), .A(n2496), .ZN(n7633) );
  OAI21_X2 U13056 ( .B1(n1569), .B2(n13245), .A(n2507), .ZN(n7634) );
  OAI21_X2 U13057 ( .B1(n1521), .B2(n13255), .A(n2416), .ZN(n7667) );
  OAI21_X2 U13058 ( .B1(n1523), .B2(n13256), .A(n2417), .ZN(n7668) );
  OAI21_X2 U13059 ( .B1(n1527), .B2(n13256), .A(n2419), .ZN(n7669) );
  OAI21_X2 U13060 ( .B1(n1529), .B2(n13256), .A(n2420), .ZN(n7670) );
  OAI21_X2 U13061 ( .B1(n1531), .B2(n13256), .A(n2421), .ZN(n7671) );
  OAI21_X2 U13062 ( .B1(n1533), .B2(n13256), .A(n2422), .ZN(n7672) );
  OAI21_X2 U13063 ( .B1(n1535), .B2(n13256), .A(n2423), .ZN(n7673) );
  OAI21_X2 U13064 ( .B1(n1537), .B2(n13256), .A(n2424), .ZN(n7674) );
  OAI21_X2 U13065 ( .B1(n1539), .B2(n13257), .A(n2425), .ZN(n7675) );
  OAI21_X2 U13066 ( .B1(n1541), .B2(n13257), .A(n2426), .ZN(n7676) );
  OAI21_X2 U13067 ( .B1(n1543), .B2(n13256), .A(n2427), .ZN(n7677) );
  OAI21_X2 U13068 ( .B1(n1545), .B2(n13257), .A(n2428), .ZN(n7678) );
  OAI21_X2 U13069 ( .B1(n1549), .B2(n13257), .A(n2430), .ZN(n7679) );
  OAI21_X2 U13070 ( .B1(n1551), .B2(n13257), .A(n2431), .ZN(n7680) );
  OAI21_X2 U13071 ( .B1(n1553), .B2(n13257), .A(n2432), .ZN(n7681) );
  OAI21_X2 U13072 ( .B1(n1555), .B2(n13257), .A(n2433), .ZN(n7682) );
  OAI21_X2 U13073 ( .B1(n1557), .B2(n13256), .A(n2434), .ZN(n7683) );
  OAI21_X2 U13074 ( .B1(n1559), .B2(n13256), .A(n2435), .ZN(n7684) );
  OAI21_X2 U13075 ( .B1(n1561), .B2(n13256), .A(n2436), .ZN(n7685) );
  OAI21_X2 U13076 ( .B1(n1563), .B2(n13255), .A(n2437), .ZN(n7686) );
  OAI21_X2 U13077 ( .B1(n1565), .B2(n13255), .A(n2438), .ZN(n7687) );
  OAI21_X2 U13078 ( .B1(n1567), .B2(n13255), .A(n2439), .ZN(n7688) );
  OAI21_X2 U13079 ( .B1(n1506), .B2(n13255), .A(n2409), .ZN(n7689) );
  OAI21_X2 U13080 ( .B1(n1509), .B2(n13255), .A(n2410), .ZN(n7690) );
  OAI21_X2 U13081 ( .B1(n1511), .B2(n13255), .A(n2411), .ZN(n7691) );
  OAI21_X2 U13082 ( .B1(n1513), .B2(n13255), .A(n2412), .ZN(n7692) );
  OAI21_X2 U13083 ( .B1(n1515), .B2(n13255), .A(n2413), .ZN(n7693) );
  OAI21_X2 U13084 ( .B1(n1517), .B2(n13255), .A(n2414), .ZN(n7694) );
  OAI21_X2 U13085 ( .B1(n1519), .B2(n13255), .A(n2415), .ZN(n7695) );
  OAI21_X2 U13086 ( .B1(n1525), .B2(n13256), .A(n2418), .ZN(n7696) );
  OAI21_X2 U13087 ( .B1(n1547), .B2(n13257), .A(n2429), .ZN(n7697) );
  OAI21_X2 U13088 ( .B1(n1569), .B2(n13255), .A(n2440), .ZN(n7698) );
  OAI21_X2 U13089 ( .B1(n1521), .B2(n13265), .A(n2348), .ZN(n7731) );
  OAI21_X2 U13090 ( .B1(n1523), .B2(n13266), .A(n2349), .ZN(n7732) );
  OAI21_X2 U13091 ( .B1(n1527), .B2(n13266), .A(n2351), .ZN(n7733) );
  OAI21_X2 U13092 ( .B1(n1529), .B2(n13266), .A(n2352), .ZN(n7734) );
  OAI21_X2 U13093 ( .B1(n1531), .B2(n13266), .A(n2353), .ZN(n7735) );
  OAI21_X2 U13094 ( .B1(n1533), .B2(n13266), .A(n2354), .ZN(n7736) );
  OAI21_X2 U13095 ( .B1(n1535), .B2(n13266), .A(n2355), .ZN(n7737) );
  OAI21_X2 U13096 ( .B1(n1537), .B2(n13266), .A(n2356), .ZN(n7738) );
  OAI21_X2 U13097 ( .B1(n1539), .B2(n13267), .A(n2357), .ZN(n7739) );
  OAI21_X2 U13098 ( .B1(n1541), .B2(n13267), .A(n2358), .ZN(n7740) );
  OAI21_X2 U13099 ( .B1(n1543), .B2(n13266), .A(n2359), .ZN(n7741) );
  OAI21_X2 U13100 ( .B1(n1545), .B2(n13267), .A(n2360), .ZN(n7742) );
  OAI21_X2 U13101 ( .B1(n1549), .B2(n13267), .A(n2362), .ZN(n7743) );
  OAI21_X2 U13102 ( .B1(n1551), .B2(n13267), .A(n2363), .ZN(n7744) );
  OAI21_X2 U13103 ( .B1(n1553), .B2(n13267), .A(n2364), .ZN(n7745) );
  OAI21_X2 U13104 ( .B1(n1555), .B2(n13267), .A(n2365), .ZN(n7746) );
  OAI21_X2 U13105 ( .B1(n1557), .B2(n13266), .A(n2366), .ZN(n7747) );
  OAI21_X2 U13106 ( .B1(n1559), .B2(n13266), .A(n2367), .ZN(n7748) );
  OAI21_X2 U13107 ( .B1(n1561), .B2(n13266), .A(n2368), .ZN(n7749) );
  OAI21_X2 U13108 ( .B1(n1563), .B2(n13265), .A(n2369), .ZN(n7750) );
  OAI21_X2 U13109 ( .B1(n1565), .B2(n13265), .A(n2370), .ZN(n7751) );
  OAI21_X2 U13110 ( .B1(n1567), .B2(n13265), .A(n2371), .ZN(n7752) );
  OAI21_X2 U13111 ( .B1(n1506), .B2(n13265), .A(n2341), .ZN(n7753) );
  OAI21_X2 U13112 ( .B1(n1509), .B2(n13265), .A(n2342), .ZN(n7754) );
  OAI21_X2 U13113 ( .B1(n1511), .B2(n13265), .A(n2343), .ZN(n7755) );
  OAI21_X2 U13114 ( .B1(n1513), .B2(n13265), .A(n2344), .ZN(n7756) );
  OAI21_X2 U13115 ( .B1(n1515), .B2(n13265), .A(n2345), .ZN(n7757) );
  OAI21_X2 U13116 ( .B1(n1517), .B2(n13265), .A(n2346), .ZN(n7758) );
  OAI21_X2 U13117 ( .B1(n1519), .B2(n13265), .A(n2347), .ZN(n7759) );
  OAI21_X2 U13118 ( .B1(n1525), .B2(n13266), .A(n2350), .ZN(n7760) );
  OAI21_X2 U13119 ( .B1(n1547), .B2(n13267), .A(n2361), .ZN(n7761) );
  OAI21_X2 U13120 ( .B1(n1569), .B2(n13265), .A(n2372), .ZN(n7762) );
  OAI21_X2 U13121 ( .B1(n13458), .B2(n13275), .A(n2282), .ZN(n7795) );
  OAI21_X2 U13122 ( .B1(n13455), .B2(n13276), .A(n2283), .ZN(n7796) );
  OAI21_X2 U13123 ( .B1(n13449), .B2(n13276), .A(n2285), .ZN(n7797) );
  OAI21_X2 U13124 ( .B1(n13446), .B2(n13276), .A(n2286), .ZN(n7798) );
  OAI21_X2 U13125 ( .B1(n13443), .B2(n13276), .A(n2287), .ZN(n7799) );
  OAI21_X2 U13126 ( .B1(n13440), .B2(n13276), .A(n2288), .ZN(n7800) );
  OAI21_X2 U13127 ( .B1(n13437), .B2(n13276), .A(n2289), .ZN(n7801) );
  OAI21_X2 U13128 ( .B1(n13434), .B2(n13276), .A(n2290), .ZN(n7802) );
  OAI21_X2 U13129 ( .B1(n13431), .B2(n13277), .A(n2291), .ZN(n7803) );
  OAI21_X2 U13130 ( .B1(n13428), .B2(n13277), .A(n2292), .ZN(n7804) );
  OAI21_X2 U13131 ( .B1(n13425), .B2(n13276), .A(n2293), .ZN(n7805) );
  OAI21_X2 U13132 ( .B1(n13422), .B2(n13277), .A(n2294), .ZN(n7806) );
  OAI21_X2 U13133 ( .B1(n13416), .B2(n13277), .A(n2296), .ZN(n7807) );
  OAI21_X2 U13134 ( .B1(n13413), .B2(n13277), .A(n2297), .ZN(n7808) );
  OAI21_X2 U13135 ( .B1(n13410), .B2(n13277), .A(n2298), .ZN(n7809) );
  OAI21_X2 U13136 ( .B1(n13407), .B2(n13277), .A(n2299), .ZN(n7810) );
  OAI21_X2 U13137 ( .B1(n13404), .B2(n13276), .A(n2300), .ZN(n7811) );
  OAI21_X2 U13138 ( .B1(n13401), .B2(n13276), .A(n2301), .ZN(n7812) );
  OAI21_X2 U13139 ( .B1(n13398), .B2(n13276), .A(n2302), .ZN(n7813) );
  OAI21_X2 U13140 ( .B1(n13395), .B2(n13275), .A(n2303), .ZN(n7814) );
  OAI21_X2 U13141 ( .B1(n13392), .B2(n13275), .A(n2304), .ZN(n7815) );
  OAI21_X2 U13142 ( .B1(n13389), .B2(n13275), .A(n2305), .ZN(n7816) );
  OAI21_X2 U13143 ( .B1(n13484), .B2(n13275), .A(n2275), .ZN(n7817) );
  OAI21_X2 U13144 ( .B1(n13476), .B2(n13275), .A(n2276), .ZN(n7818) );
  OAI21_X2 U13145 ( .B1(n13473), .B2(n13275), .A(n2277), .ZN(n7819) );
  OAI21_X2 U13146 ( .B1(n13470), .B2(n13275), .A(n2278), .ZN(n7820) );
  OAI21_X2 U13147 ( .B1(n13467), .B2(n13275), .A(n2279), .ZN(n7821) );
  OAI21_X2 U13148 ( .B1(n13464), .B2(n13275), .A(n2280), .ZN(n7822) );
  OAI21_X2 U13149 ( .B1(n13461), .B2(n13275), .A(n2281), .ZN(n7823) );
  OAI21_X2 U13150 ( .B1(n13452), .B2(n13276), .A(n2284), .ZN(n7824) );
  OAI21_X2 U13151 ( .B1(n13419), .B2(n13277), .A(n2295), .ZN(n7825) );
  OAI21_X2 U13152 ( .B1(n13386), .B2(n13275), .A(n2306), .ZN(n7826) );
  OAI21_X2 U13153 ( .B1(n13458), .B2(n13290), .A(n2181), .ZN(n7859) );
  OAI21_X2 U13154 ( .B1(n13455), .B2(n13291), .A(n2182), .ZN(n7860) );
  OAI21_X2 U13155 ( .B1(n13449), .B2(n13291), .A(n2184), .ZN(n7861) );
  OAI21_X2 U13156 ( .B1(n13446), .B2(n13291), .A(n2185), .ZN(n7862) );
  OAI21_X2 U13157 ( .B1(n13443), .B2(n13291), .A(n2186), .ZN(n7863) );
  OAI21_X2 U13158 ( .B1(n13440), .B2(n13291), .A(n2187), .ZN(n7864) );
  OAI21_X2 U13159 ( .B1(n13437), .B2(n13291), .A(n2188), .ZN(n7865) );
  OAI21_X2 U13160 ( .B1(n13434), .B2(n13291), .A(n2189), .ZN(n7866) );
  OAI21_X2 U13161 ( .B1(n13431), .B2(n13292), .A(n2190), .ZN(n7867) );
  OAI21_X2 U13162 ( .B1(n13428), .B2(n13292), .A(n2191), .ZN(n7868) );
  OAI21_X2 U13163 ( .B1(n13425), .B2(n13291), .A(n2192), .ZN(n7869) );
  OAI21_X2 U13164 ( .B1(n13422), .B2(n13292), .A(n2193), .ZN(n7870) );
  OAI21_X2 U13165 ( .B1(n13416), .B2(n13292), .A(n2195), .ZN(n7871) );
  OAI21_X2 U13166 ( .B1(n13413), .B2(n13292), .A(n2196), .ZN(n7872) );
  OAI21_X2 U13167 ( .B1(n13410), .B2(n13292), .A(n2197), .ZN(n7873) );
  OAI21_X2 U13168 ( .B1(n13407), .B2(n13292), .A(n2198), .ZN(n7874) );
  OAI21_X2 U13169 ( .B1(n13404), .B2(n13291), .A(n2199), .ZN(n7875) );
  OAI21_X2 U13170 ( .B1(n13401), .B2(n13291), .A(n2200), .ZN(n7876) );
  OAI21_X2 U13171 ( .B1(n13398), .B2(n13291), .A(n2201), .ZN(n7877) );
  OAI21_X2 U13172 ( .B1(n13395), .B2(n13290), .A(n2202), .ZN(n7878) );
  OAI21_X2 U13173 ( .B1(n13392), .B2(n13290), .A(n2203), .ZN(n7879) );
  OAI21_X2 U13174 ( .B1(n13389), .B2(n13290), .A(n2204), .ZN(n7880) );
  OAI21_X2 U13175 ( .B1(n13484), .B2(n13290), .A(n2174), .ZN(n7881) );
  OAI21_X2 U13176 ( .B1(n13476), .B2(n13290), .A(n2175), .ZN(n7882) );
  OAI21_X2 U13177 ( .B1(n13473), .B2(n13290), .A(n2176), .ZN(n7883) );
  OAI21_X2 U13178 ( .B1(n13470), .B2(n13290), .A(n2177), .ZN(n7884) );
  OAI21_X2 U13179 ( .B1(n13467), .B2(n13290), .A(n2178), .ZN(n7885) );
  OAI21_X2 U13180 ( .B1(n13464), .B2(n13290), .A(n2179), .ZN(n7886) );
  OAI21_X2 U13181 ( .B1(n13461), .B2(n13290), .A(n2180), .ZN(n7887) );
  OAI21_X2 U13182 ( .B1(n13452), .B2(n13291), .A(n2183), .ZN(n7888) );
  OAI21_X2 U13183 ( .B1(n13419), .B2(n13292), .A(n2194), .ZN(n7889) );
  OAI21_X2 U13184 ( .B1(n13386), .B2(n13290), .A(n2205), .ZN(n7890) );
  OAI21_X2 U13185 ( .B1(n13458), .B2(n13300), .A(n2115), .ZN(n7923) );
  OAI21_X2 U13186 ( .B1(n13455), .B2(n13301), .A(n2116), .ZN(n7924) );
  OAI21_X2 U13187 ( .B1(n13449), .B2(n13301), .A(n2118), .ZN(n7925) );
  OAI21_X2 U13188 ( .B1(n13446), .B2(n13301), .A(n2119), .ZN(n7926) );
  OAI21_X2 U13189 ( .B1(n13443), .B2(n13301), .A(n2120), .ZN(n7927) );
  OAI21_X2 U13190 ( .B1(n13440), .B2(n13301), .A(n2121), .ZN(n7928) );
  OAI21_X2 U13191 ( .B1(n13437), .B2(n13301), .A(n2122), .ZN(n7929) );
  OAI21_X2 U13192 ( .B1(n13434), .B2(n13301), .A(n2123), .ZN(n7930) );
  OAI21_X2 U13193 ( .B1(n13431), .B2(n13302), .A(n2124), .ZN(n7931) );
  OAI21_X2 U13194 ( .B1(n13428), .B2(n13302), .A(n2125), .ZN(n7932) );
  OAI21_X2 U13195 ( .B1(n13425), .B2(n13301), .A(n2126), .ZN(n7933) );
  OAI21_X2 U13196 ( .B1(n13422), .B2(n13302), .A(n2127), .ZN(n7934) );
  OAI21_X2 U13197 ( .B1(n13416), .B2(n13302), .A(n2129), .ZN(n7935) );
  OAI21_X2 U13198 ( .B1(n13413), .B2(n13302), .A(n2130), .ZN(n7936) );
  OAI21_X2 U13199 ( .B1(n13410), .B2(n13302), .A(n2131), .ZN(n7937) );
  OAI21_X2 U13200 ( .B1(n13407), .B2(n13302), .A(n2132), .ZN(n7938) );
  OAI21_X2 U13201 ( .B1(n13404), .B2(n13301), .A(n2133), .ZN(n7939) );
  OAI21_X2 U13202 ( .B1(n13401), .B2(n13301), .A(n2134), .ZN(n7940) );
  OAI21_X2 U13203 ( .B1(n13398), .B2(n13301), .A(n2135), .ZN(n7941) );
  OAI21_X2 U13204 ( .B1(n13395), .B2(n13300), .A(n2136), .ZN(n7942) );
  OAI21_X2 U13205 ( .B1(n13392), .B2(n13300), .A(n2137), .ZN(n7943) );
  OAI21_X2 U13206 ( .B1(n13389), .B2(n13300), .A(n2138), .ZN(n7944) );
  OAI21_X2 U13207 ( .B1(n13484), .B2(n13300), .A(n2108), .ZN(n7945) );
  OAI21_X2 U13208 ( .B1(n13476), .B2(n13300), .A(n2109), .ZN(n7946) );
  OAI21_X2 U13209 ( .B1(n13473), .B2(n13300), .A(n2110), .ZN(n7947) );
  OAI21_X2 U13210 ( .B1(n13470), .B2(n13300), .A(n2111), .ZN(n7948) );
  OAI21_X2 U13211 ( .B1(n13467), .B2(n13300), .A(n2112), .ZN(n7949) );
  OAI21_X2 U13212 ( .B1(n13464), .B2(n13300), .A(n2113), .ZN(n7950) );
  OAI21_X2 U13213 ( .B1(n13461), .B2(n13300), .A(n2114), .ZN(n7951) );
  OAI21_X2 U13214 ( .B1(n13452), .B2(n13301), .A(n2117), .ZN(n7952) );
  OAI21_X2 U13215 ( .B1(n13419), .B2(n13302), .A(n2128), .ZN(n7953) );
  OAI21_X2 U13216 ( .B1(n13386), .B2(n13300), .A(n2139), .ZN(n7954) );
  OAI21_X2 U13217 ( .B1(n13458), .B2(n13310), .A(n2048), .ZN(n7987) );
  OAI21_X2 U13218 ( .B1(n13455), .B2(n13311), .A(n2049), .ZN(n7988) );
  OAI21_X2 U13219 ( .B1(n13449), .B2(n13311), .A(n2051), .ZN(n7989) );
  OAI21_X2 U13220 ( .B1(n13446), .B2(n13311), .A(n2052), .ZN(n7990) );
  OAI21_X2 U13221 ( .B1(n13443), .B2(n13311), .A(n2053), .ZN(n7991) );
  OAI21_X2 U13222 ( .B1(n13440), .B2(n13311), .A(n2054), .ZN(n7992) );
  OAI21_X2 U13223 ( .B1(n13437), .B2(n13311), .A(n2055), .ZN(n7993) );
  OAI21_X2 U13224 ( .B1(n13434), .B2(n13311), .A(n2056), .ZN(n7994) );
  OAI21_X2 U13225 ( .B1(n13431), .B2(n13312), .A(n2057), .ZN(n7995) );
  OAI21_X2 U13226 ( .B1(n13428), .B2(n13312), .A(n2058), .ZN(n7996) );
  OAI21_X2 U13227 ( .B1(n13425), .B2(n13311), .A(n2059), .ZN(n7997) );
  OAI21_X2 U13228 ( .B1(n13422), .B2(n13312), .A(n2060), .ZN(n7998) );
  OAI21_X2 U13229 ( .B1(n13416), .B2(n13312), .A(n2062), .ZN(n7999) );
  OAI21_X2 U13230 ( .B1(n13413), .B2(n13312), .A(n2063), .ZN(n8000) );
  OAI21_X2 U13231 ( .B1(n13410), .B2(n13312), .A(n2064), .ZN(n8001) );
  OAI21_X2 U13232 ( .B1(n13407), .B2(n13312), .A(n2065), .ZN(n8002) );
  OAI21_X2 U13233 ( .B1(n13404), .B2(n13311), .A(n2066), .ZN(n8003) );
  OAI21_X2 U13234 ( .B1(n13401), .B2(n13311), .A(n2067), .ZN(n8004) );
  OAI21_X2 U13235 ( .B1(n13398), .B2(n13311), .A(n2068), .ZN(n8005) );
  OAI21_X2 U13236 ( .B1(n13395), .B2(n13310), .A(n2069), .ZN(n8006) );
  OAI21_X2 U13237 ( .B1(n13392), .B2(n13310), .A(n2070), .ZN(n8007) );
  OAI21_X2 U13238 ( .B1(n13389), .B2(n13310), .A(n2071), .ZN(n8008) );
  OAI21_X2 U13239 ( .B1(n13484), .B2(n13310), .A(n2041), .ZN(n8009) );
  OAI21_X2 U13240 ( .B1(n13476), .B2(n13310), .A(n2042), .ZN(n8010) );
  OAI21_X2 U13241 ( .B1(n13473), .B2(n13310), .A(n2043), .ZN(n8011) );
  OAI21_X2 U13242 ( .B1(n13470), .B2(n13310), .A(n2044), .ZN(n8012) );
  OAI21_X2 U13243 ( .B1(n13467), .B2(n13310), .A(n2045), .ZN(n8013) );
  OAI21_X2 U13244 ( .B1(n13464), .B2(n13310), .A(n2046), .ZN(n8014) );
  OAI21_X2 U13245 ( .B1(n13461), .B2(n13310), .A(n2047), .ZN(n8015) );
  OAI21_X2 U13246 ( .B1(n13452), .B2(n13311), .A(n2050), .ZN(n8016) );
  OAI21_X2 U13247 ( .B1(n13419), .B2(n13312), .A(n2061), .ZN(n8017) );
  OAI21_X2 U13248 ( .B1(n13386), .B2(n13310), .A(n2072), .ZN(n8018) );
  OAI21_X2 U13249 ( .B1(n13458), .B2(n13320), .A(n1982), .ZN(n8051) );
  OAI21_X2 U13250 ( .B1(n13455), .B2(n13321), .A(n1983), .ZN(n8052) );
  OAI21_X2 U13251 ( .B1(n13449), .B2(n13321), .A(n1985), .ZN(n8053) );
  OAI21_X2 U13252 ( .B1(n13446), .B2(n13321), .A(n1986), .ZN(n8054) );
  OAI21_X2 U13253 ( .B1(n13443), .B2(n13321), .A(n1987), .ZN(n8055) );
  OAI21_X2 U13254 ( .B1(n13440), .B2(n13321), .A(n1988), .ZN(n8056) );
  OAI21_X2 U13255 ( .B1(n13437), .B2(n13321), .A(n1989), .ZN(n8057) );
  OAI21_X2 U13256 ( .B1(n13434), .B2(n13321), .A(n1990), .ZN(n8058) );
  OAI21_X2 U13257 ( .B1(n13431), .B2(n13322), .A(n1991), .ZN(n8059) );
  OAI21_X2 U13258 ( .B1(n13428), .B2(n13322), .A(n1992), .ZN(n8060) );
  OAI21_X2 U13259 ( .B1(n13425), .B2(n13321), .A(n1993), .ZN(n8061) );
  OAI21_X2 U13260 ( .B1(n13422), .B2(n13322), .A(n1994), .ZN(n8062) );
  OAI21_X2 U13261 ( .B1(n13416), .B2(n13322), .A(n1996), .ZN(n8063) );
  OAI21_X2 U13262 ( .B1(n13413), .B2(n13322), .A(n1997), .ZN(n8064) );
  OAI21_X2 U13263 ( .B1(n13410), .B2(n13322), .A(n1998), .ZN(n8065) );
  OAI21_X2 U13264 ( .B1(n13407), .B2(n13322), .A(n1999), .ZN(n8066) );
  OAI21_X2 U13265 ( .B1(n13404), .B2(n13321), .A(n2000), .ZN(n8067) );
  OAI21_X2 U13266 ( .B1(n13401), .B2(n13321), .A(n2001), .ZN(n8068) );
  OAI21_X2 U13267 ( .B1(n13398), .B2(n13321), .A(n2002), .ZN(n8069) );
  OAI21_X2 U13268 ( .B1(n13395), .B2(n13320), .A(n2003), .ZN(n8070) );
  OAI21_X2 U13269 ( .B1(n13392), .B2(n13320), .A(n2004), .ZN(n8071) );
  OAI21_X2 U13270 ( .B1(n13389), .B2(n13320), .A(n2005), .ZN(n8072) );
  OAI21_X2 U13271 ( .B1(n13484), .B2(n13320), .A(n1975), .ZN(n8073) );
  OAI21_X2 U13272 ( .B1(n13476), .B2(n13320), .A(n1976), .ZN(n8074) );
  OAI21_X2 U13273 ( .B1(n13473), .B2(n13320), .A(n1977), .ZN(n8075) );
  OAI21_X2 U13274 ( .B1(n13470), .B2(n13320), .A(n1978), .ZN(n8076) );
  OAI21_X2 U13275 ( .B1(n13467), .B2(n13320), .A(n1979), .ZN(n8077) );
  OAI21_X2 U13276 ( .B1(n13464), .B2(n13320), .A(n1980), .ZN(n8078) );
  OAI21_X2 U13277 ( .B1(n13461), .B2(n13320), .A(n1981), .ZN(n8079) );
  OAI21_X2 U13278 ( .B1(n13452), .B2(n13321), .A(n1984), .ZN(n8080) );
  OAI21_X2 U13279 ( .B1(n13419), .B2(n13322), .A(n1995), .ZN(n8081) );
  OAI21_X2 U13280 ( .B1(n13386), .B2(n13320), .A(n2006), .ZN(n8082) );
  OAI21_X2 U13281 ( .B1(n13457), .B2(n13330), .A(n1914), .ZN(n8115) );
  OAI21_X2 U13282 ( .B1(n13454), .B2(n13331), .A(n1915), .ZN(n8116) );
  OAI21_X2 U13283 ( .B1(n13448), .B2(n13331), .A(n1917), .ZN(n8117) );
  OAI21_X2 U13284 ( .B1(n13445), .B2(n13331), .A(n1918), .ZN(n8118) );
  OAI21_X2 U13285 ( .B1(n13442), .B2(n13331), .A(n1919), .ZN(n8119) );
  OAI21_X2 U13286 ( .B1(n13439), .B2(n13331), .A(n1920), .ZN(n8120) );
  OAI21_X2 U13287 ( .B1(n13436), .B2(n13331), .A(n1921), .ZN(n8121) );
  OAI21_X2 U13288 ( .B1(n13433), .B2(n13331), .A(n1922), .ZN(n8122) );
  OAI21_X2 U13289 ( .B1(n13430), .B2(n13332), .A(n1923), .ZN(n8123) );
  OAI21_X2 U13290 ( .B1(n13427), .B2(n13332), .A(n1924), .ZN(n8124) );
  OAI21_X2 U13291 ( .B1(n13424), .B2(n13331), .A(n1925), .ZN(n8125) );
  OAI21_X2 U13292 ( .B1(n13421), .B2(n13332), .A(n1926), .ZN(n8126) );
  OAI21_X2 U13293 ( .B1(n13415), .B2(n13332), .A(n1928), .ZN(n8127) );
  OAI21_X2 U13294 ( .B1(n13412), .B2(n13332), .A(n1929), .ZN(n8128) );
  OAI21_X2 U13295 ( .B1(n13409), .B2(n13332), .A(n1930), .ZN(n8129) );
  OAI21_X2 U13296 ( .B1(n13406), .B2(n13332), .A(n1931), .ZN(n8130) );
  OAI21_X2 U13297 ( .B1(n13403), .B2(n13331), .A(n1932), .ZN(n8131) );
  OAI21_X2 U13298 ( .B1(n13400), .B2(n13331), .A(n1933), .ZN(n8132) );
  OAI21_X2 U13299 ( .B1(n13397), .B2(n13331), .A(n1934), .ZN(n8133) );
  OAI21_X2 U13300 ( .B1(n13394), .B2(n13330), .A(n1935), .ZN(n8134) );
  OAI21_X2 U13301 ( .B1(n13391), .B2(n13330), .A(n1936), .ZN(n8135) );
  OAI21_X2 U13302 ( .B1(n13388), .B2(n13330), .A(n1937), .ZN(n8136) );
  OAI21_X2 U13303 ( .B1(n13483), .B2(n13330), .A(n1907), .ZN(n8137) );
  OAI21_X2 U13304 ( .B1(n13475), .B2(n13330), .A(n1908), .ZN(n8138) );
  OAI21_X2 U13305 ( .B1(n13472), .B2(n13330), .A(n1909), .ZN(n8139) );
  OAI21_X2 U13306 ( .B1(n13469), .B2(n13330), .A(n1910), .ZN(n8140) );
  OAI21_X2 U13307 ( .B1(n13466), .B2(n13330), .A(n1911), .ZN(n8141) );
  OAI21_X2 U13308 ( .B1(n13463), .B2(n13330), .A(n1912), .ZN(n8142) );
  OAI21_X2 U13309 ( .B1(n13460), .B2(n13330), .A(n1913), .ZN(n8143) );
  OAI21_X2 U13310 ( .B1(n13451), .B2(n13331), .A(n1916), .ZN(n8144) );
  OAI21_X2 U13311 ( .B1(n13418), .B2(n13332), .A(n1927), .ZN(n8145) );
  OAI21_X2 U13312 ( .B1(n13385), .B2(n13330), .A(n1938), .ZN(n8146) );
  OAI21_X2 U13313 ( .B1(n13457), .B2(n13345), .A(n1815), .ZN(n8179) );
  OAI21_X2 U13314 ( .B1(n13454), .B2(n13346), .A(n1816), .ZN(n8180) );
  OAI21_X2 U13315 ( .B1(n13448), .B2(n13346), .A(n1818), .ZN(n8181) );
  OAI21_X2 U13316 ( .B1(n13445), .B2(n13346), .A(n1819), .ZN(n8182) );
  OAI21_X2 U13317 ( .B1(n13442), .B2(n13346), .A(n1820), .ZN(n8183) );
  OAI21_X2 U13318 ( .B1(n13439), .B2(n13346), .A(n1821), .ZN(n8184) );
  OAI21_X2 U13319 ( .B1(n13436), .B2(n13346), .A(n1822), .ZN(n8185) );
  OAI21_X2 U13320 ( .B1(n13433), .B2(n13346), .A(n1823), .ZN(n8186) );
  OAI21_X2 U13321 ( .B1(n13430), .B2(n13347), .A(n1824), .ZN(n8187) );
  OAI21_X2 U13322 ( .B1(n13427), .B2(n13347), .A(n1825), .ZN(n8188) );
  OAI21_X2 U13323 ( .B1(n13424), .B2(n13346), .A(n1826), .ZN(n8189) );
  OAI21_X2 U13324 ( .B1(n13421), .B2(n13347), .A(n1827), .ZN(n8190) );
  OAI21_X2 U13325 ( .B1(n13415), .B2(n13347), .A(n1829), .ZN(n8191) );
  OAI21_X2 U13326 ( .B1(n13412), .B2(n13347), .A(n1830), .ZN(n8192) );
  OAI21_X2 U13327 ( .B1(n13409), .B2(n13347), .A(n1831), .ZN(n8193) );
  OAI21_X2 U13328 ( .B1(n13406), .B2(n13347), .A(n1832), .ZN(n8194) );
  OAI21_X2 U13329 ( .B1(n13403), .B2(n13346), .A(n1833), .ZN(n8195) );
  OAI21_X2 U13330 ( .B1(n13400), .B2(n13346), .A(n1834), .ZN(n8196) );
  OAI21_X2 U13331 ( .B1(n13397), .B2(n13346), .A(n1835), .ZN(n8197) );
  OAI21_X2 U13332 ( .B1(n13394), .B2(n13345), .A(n1836), .ZN(n8198) );
  OAI21_X2 U13333 ( .B1(n13391), .B2(n13345), .A(n1837), .ZN(n8199) );
  OAI21_X2 U13334 ( .B1(n13388), .B2(n13345), .A(n1838), .ZN(n8200) );
  OAI21_X2 U13335 ( .B1(n13483), .B2(n13345), .A(n1808), .ZN(n8201) );
  OAI21_X2 U13336 ( .B1(n13475), .B2(n13345), .A(n1809), .ZN(n8202) );
  OAI21_X2 U13337 ( .B1(n13472), .B2(n13345), .A(n1810), .ZN(n8203) );
  OAI21_X2 U13338 ( .B1(n13469), .B2(n13345), .A(n1811), .ZN(n8204) );
  OAI21_X2 U13339 ( .B1(n13466), .B2(n13345), .A(n1812), .ZN(n8205) );
  OAI21_X2 U13340 ( .B1(n13463), .B2(n13345), .A(n1813), .ZN(n8206) );
  OAI21_X2 U13341 ( .B1(n13460), .B2(n13345), .A(n1814), .ZN(n8207) );
  OAI21_X2 U13342 ( .B1(n13451), .B2(n13346), .A(n1817), .ZN(n8208) );
  OAI21_X2 U13343 ( .B1(n13418), .B2(n13347), .A(n1828), .ZN(n8209) );
  OAI21_X2 U13344 ( .B1(n13385), .B2(n13345), .A(n1839), .ZN(n8210) );
  MUX2_X2 U13345 ( .A(decode_regfile_intregs_31__0_), .B(
        decode_regfile_intregs_30__0_), .S(n13802), .Z(n8826) );
  MUX2_X2 U13346 ( .A(decode_regfile_intregs_31__0_), .B(
        decode_regfile_intregs_30__0_), .S(n8810), .Z(n10961) );
  OAI22_X2 U13347 ( .A1(execstage_Imm32[24]), .A2(n13787), .B1(n13788), .B2(
        busB_1[24]), .ZN(n3480) );
  AND4_X2 U13348 ( .A1(execstage_AluCtrl[0]), .A2(n8720), .A3(n8697), .A4(
        n8660), .ZN(n8818) );
  AOI21_X2 U13349 ( .B1(n6085), .B2(n6164), .A(n6165), .ZN(n6163) );
  NOR3_X2 U13350 ( .A1(n3442), .A2(n16426), .A3(n8735), .ZN(n6165) );
  NAND3_X2 U13351 ( .A1(n4100), .A2(n4101), .A3(n4102), .ZN(n3236) );
  NAND3_X2 U13352 ( .A1(n4389), .A2(n4390), .A3(n4391), .ZN(n3647) );
  AOI21_X2 U13353 ( .B1(execstage_AluCtrl[0]), .B2(n6056), .A(n6057), .ZN(
        n6055) );
  NAND3_X2 U13354 ( .A1(n13129), .A2(execstage_ALU_ra_row2_31_), .A3(n13197), 
        .ZN(n6178) );
  OAI21_X2 U13355 ( .B1(execstage_BusA[27]), .B2(n3209), .A(n6088), .ZN(n6086)
         );
  NOR3_X2 U13356 ( .A1(execstage_AluCtrl[2]), .A2(execstage_AluCtrl[3]), .A3(
        execstage_AluCtrl[0]), .ZN(n6045) );
  NOR3_X2 U13357 ( .A1(execstage_AluCtrl[0]), .A2(execstage_AluCtrl[1]), .A3(
        n8697), .ZN(n6051) );
  NOR2_X2 U13358 ( .A1(n6056), .A2(execstage_AluCtrl[0]), .ZN(n6057) );
  NOR3_X2 U13359 ( .A1(n3442), .A2(execstage_BusA[28]), .A3(n3455), .ZN(n6087)
         );
  OAI21_X2 U13360 ( .B1(n13804), .B2(n134), .A(n135), .ZN(
        execstage_register_N6) );
  AOI222_X1 U13361 ( .A1(n16602), .A2(n137), .B1(n138), .B2(n139), .C1(n16598), 
        .C2(n141), .ZN(n134) );
  NOR2_X2 U13362 ( .A1(n8754), .A2(rw_3[1]), .ZN(n800) );
  NOR2_X2 U13363 ( .A1(rw_3[1]), .A2(rw_3[0]), .ZN(n834) );
  NOR2_X2 U13364 ( .A1(imm32_0[9]), .A2(imm32_0[8]), .ZN(n2677) );
  NOR2_X2 U13365 ( .A1(rw_3[3]), .A2(rw_3[2]), .ZN(n664) );
  NOR2_X2 U13366 ( .A1(n8729), .A2(rw_3[3]), .ZN(n530) );
  NOR2_X2 U13367 ( .A1(n8752), .A2(rw_3[2]), .ZN(n461) );
  NOR2_X2 U13368 ( .A1(n8726), .A2(imm32_0[0]), .ZN(n2657) );
  OAI21_X2 U13369 ( .B1(n13488), .B2(n13486), .A(wrenable), .ZN(n1270) );
  OAI21_X2 U13370 ( .B1(n13228), .B2(n16357), .A(wrenable), .ZN(n2373) );
  OAI21_X2 U13371 ( .B1(instruction_2[28]), .B2(n8762), .A(instruction_2[27]), 
        .ZN(n6193) );
  AOI21_X2 U13372 ( .B1(n6189), .B2(n6190), .A(instruction_2[30]), .ZN(N139)
         );
  NAND3_X2 U13373 ( .A1(n6193), .A2(n8797), .A3(instruction_2[31]), .ZN(n6189)
         );
  NOR2_X2 U13374 ( .A1(n1270), .A2(rw_3[4]), .ZN(n1370) );
  NOR2_X2 U13375 ( .A1(n2373), .A2(rw_3[4]), .ZN(n1738) );
  NOR2_X2 U13376 ( .A1(instruction_2[31]), .A2(n8762), .ZN(n6191) );
  NAND2_X2 U13377 ( .A1(fpoint_3[1]), .A2(fpoint_3[0]), .ZN(n8819) );
  OR2_X2 U13378 ( .A1(fpoint_3[0]), .A2(fpoint_3[1]), .ZN(n8820) );
  OR2_X2 U13379 ( .A1(n8724), .A2(fpoint_3[0]), .ZN(n8821) );
  NOR3_X2 U13380 ( .A1(imm32_0[4]), .A2(imm32_0[5]), .A3(n147), .ZN(n2656) );
  AOI211_X2 U13381 ( .C1(n138), .C2(n2643), .A(n306), .B(n16601), .ZN(n2642)
         );
  NAND3_X2 U13382 ( .A1(imm32_0[3]), .A2(n8727), .A3(n16587), .ZN(n2647) );
  NOR2_X2 U13383 ( .A1(fwdB[0]), .A2(n13804), .ZN(n266) );
  NAND3_X2 U13384 ( .A1(imm32_0[3]), .A2(imm32_0[2]), .A3(n16587), .ZN(n2645)
         );
  NAND3_X2 U13385 ( .A1(n2657), .A2(imm32_0[2]), .A3(n2674), .ZN(n2652) );
  AOI21_X2 U13386 ( .B1(imm32_0[3]), .B2(imm32_0[4]), .A(imm32_0[5]), .ZN(
        n2674) );
  NOR2_X2 U13387 ( .A1(fwdA[0]), .A2(fwdA[1]), .ZN(n393) );
  AND2_X2 U13388 ( .A1(fwdA[1]), .A2(n16217), .ZN(n8822) );
  AND2_X2 U13389 ( .A1(fwdB[1]), .A2(n266), .ZN(n8823) );
  NOR2_X2 U13390 ( .A1(n16217), .A2(fwdA[1]), .ZN(n8824) );
  AND3_X2 U13391 ( .A1(n16547), .A2(n13809), .A3(fwdB[0]), .ZN(n8825) );
  INV_X4 U13392 ( .A(stall), .ZN(n13803) );
  NAND3_X2 U13393 ( .A1(n2665), .A2(n8726), .A3(imm32_0[0]), .ZN(n2673) );
  OAI21_X2 U13394 ( .B1(N15), .B2(n16371), .A(n16214), .ZN(N46) );
  MUX2_X2 U13395 ( .A(decode_regfile_intregs_28__0_), .B(
        decode_regfile_intregs_29__0_), .S(n10777), .Z(n8827) );
  MUX2_X2 U13396 ( .A(n8827), .B(n8826), .S(n10879), .Z(n8828) );
  MUX2_X2 U13397 ( .A(decode_regfile_intregs_26__0_), .B(
        decode_regfile_intregs_27__0_), .S(n10777), .Z(n8829) );
  MUX2_X2 U13398 ( .A(decode_regfile_intregs_24__0_), .B(
        decode_regfile_intregs_25__0_), .S(n10777), .Z(n8830) );
  MUX2_X2 U13399 ( .A(n8830), .B(n8829), .S(n10879), .Z(n8831) );
  MUX2_X2 U13400 ( .A(n8831), .B(n8828), .S(n10921), .Z(n8832) );
  MUX2_X2 U13401 ( .A(decode_regfile_intregs_22__0_), .B(
        decode_regfile_intregs_23__0_), .S(n10777), .Z(n8833) );
  MUX2_X2 U13402 ( .A(decode_regfile_intregs_20__0_), .B(
        decode_regfile_intregs_21__0_), .S(n10777), .Z(n8834) );
  MUX2_X2 U13403 ( .A(n8834), .B(n8833), .S(n10879), .Z(n8835) );
  MUX2_X2 U13404 ( .A(decode_regfile_intregs_18__0_), .B(
        decode_regfile_intregs_19__0_), .S(n10777), .Z(n8836) );
  MUX2_X2 U13405 ( .A(decode_regfile_intregs_16__0_), .B(
        decode_regfile_intregs_17__0_), .S(n10777), .Z(n8837) );
  MUX2_X2 U13406 ( .A(n8837), .B(n8836), .S(n10879), .Z(n8838) );
  MUX2_X2 U13407 ( .A(n8838), .B(n8835), .S(n10921), .Z(n8839) );
  MUX2_X2 U13408 ( .A(n8839), .B(n8832), .S(decode_rs2_3_), .Z(n8840) );
  MUX2_X2 U13409 ( .A(decode_regfile_intregs_14__0_), .B(
        decode_regfile_intregs_15__0_), .S(n10777), .Z(n8841) );
  MUX2_X2 U13410 ( .A(decode_regfile_intregs_12__0_), .B(
        decode_regfile_intregs_13__0_), .S(n10777), .Z(n8842) );
  MUX2_X2 U13411 ( .A(n8842), .B(n8841), .S(n10879), .Z(n8843) );
  MUX2_X2 U13412 ( .A(decode_regfile_intregs_10__0_), .B(
        decode_regfile_intregs_11__0_), .S(n10777), .Z(n8844) );
  MUX2_X2 U13413 ( .A(decode_regfile_intregs_8__0_), .B(
        decode_regfile_intregs_9__0_), .S(n10777), .Z(n8845) );
  MUX2_X2 U13414 ( .A(n8845), .B(n8844), .S(n10879), .Z(n8846) );
  MUX2_X2 U13415 ( .A(n8846), .B(n8843), .S(n10921), .Z(n8847) );
  MUX2_X2 U13416 ( .A(decode_regfile_intregs_6__0_), .B(
        decode_regfile_intregs_7__0_), .S(n10778), .Z(n8848) );
  MUX2_X2 U13417 ( .A(decode_regfile_intregs_4__0_), .B(
        decode_regfile_intregs_5__0_), .S(n10778), .Z(n8849) );
  MUX2_X2 U13418 ( .A(n8849), .B(n8848), .S(n10880), .Z(n8850) );
  MUX2_X2 U13419 ( .A(decode_regfile_intregs_2__0_), .B(
        decode_regfile_intregs_3__0_), .S(n10778), .Z(n8851) );
  MUX2_X2 U13420 ( .A(decode_regfile_intregs_0__0_), .B(
        decode_regfile_intregs_1__0_), .S(n10778), .Z(n8852) );
  MUX2_X2 U13421 ( .A(n8852), .B(n8851), .S(n10880), .Z(n8853) );
  MUX2_X2 U13422 ( .A(n8853), .B(n8850), .S(n10922), .Z(n8854) );
  MUX2_X2 U13423 ( .A(n8854), .B(n8847), .S(decode_rs2_3_), .Z(n8855) );
  MUX2_X2 U13424 ( .A(n8855), .B(n8840), .S(decode_rs2_4_), .Z(
        decode_regfile_N91) );
  MUX2_X2 U13425 ( .A(decode_regfile_intregs_30__1_), .B(
        decode_regfile_intregs_31__1_), .S(n10778), .Z(n8856) );
  MUX2_X2 U13426 ( .A(decode_regfile_intregs_28__1_), .B(
        decode_regfile_intregs_29__1_), .S(n10778), .Z(n8857) );
  MUX2_X2 U13427 ( .A(n8857), .B(n8856), .S(n10880), .Z(n8858) );
  MUX2_X2 U13428 ( .A(decode_regfile_intregs_26__1_), .B(
        decode_regfile_intregs_27__1_), .S(n10778), .Z(n8859) );
  MUX2_X2 U13429 ( .A(decode_regfile_intregs_24__1_), .B(
        decode_regfile_intregs_25__1_), .S(n10778), .Z(n8860) );
  MUX2_X2 U13430 ( .A(n8860), .B(n8859), .S(n10880), .Z(n8861) );
  MUX2_X2 U13431 ( .A(n8861), .B(n8858), .S(n10922), .Z(n8862) );
  MUX2_X2 U13432 ( .A(decode_regfile_intregs_22__1_), .B(
        decode_regfile_intregs_23__1_), .S(n10778), .Z(n8863) );
  MUX2_X2 U13433 ( .A(decode_regfile_intregs_20__1_), .B(
        decode_regfile_intregs_21__1_), .S(n10778), .Z(n8864) );
  MUX2_X2 U13434 ( .A(n8864), .B(n8863), .S(n10880), .Z(n8865) );
  MUX2_X2 U13435 ( .A(decode_regfile_intregs_18__1_), .B(
        decode_regfile_intregs_19__1_), .S(n10778), .Z(n8866) );
  MUX2_X2 U13436 ( .A(decode_regfile_intregs_16__1_), .B(
        decode_regfile_intregs_17__1_), .S(n10779), .Z(n8867) );
  MUX2_X2 U13437 ( .A(n8867), .B(n8866), .S(n10880), .Z(n8868) );
  MUX2_X2 U13438 ( .A(n8868), .B(n8865), .S(n10922), .Z(n8869) );
  MUX2_X2 U13439 ( .A(n8869), .B(n8862), .S(decode_rs2_3_), .Z(n8870) );
  MUX2_X2 U13440 ( .A(decode_regfile_intregs_14__1_), .B(
        decode_regfile_intregs_15__1_), .S(n10779), .Z(n8871) );
  MUX2_X2 U13441 ( .A(decode_regfile_intregs_12__1_), .B(
        decode_regfile_intregs_13__1_), .S(n10779), .Z(n8872) );
  MUX2_X2 U13442 ( .A(n8872), .B(n8871), .S(n10880), .Z(n8873) );
  MUX2_X2 U13443 ( .A(decode_regfile_intregs_10__1_), .B(
        decode_regfile_intregs_11__1_), .S(n10779), .Z(n8874) );
  MUX2_X2 U13444 ( .A(decode_regfile_intregs_8__1_), .B(
        decode_regfile_intregs_9__1_), .S(n10779), .Z(n8875) );
  MUX2_X2 U13445 ( .A(n8875), .B(n8874), .S(n10880), .Z(n8876) );
  MUX2_X2 U13446 ( .A(n8876), .B(n8873), .S(n10922), .Z(n8877) );
  MUX2_X2 U13447 ( .A(decode_regfile_intregs_6__1_), .B(
        decode_regfile_intregs_7__1_), .S(n10779), .Z(n8878) );
  MUX2_X2 U13448 ( .A(decode_regfile_intregs_4__1_), .B(
        decode_regfile_intregs_5__1_), .S(n10779), .Z(n8879) );
  MUX2_X2 U13449 ( .A(n8879), .B(n8878), .S(n10880), .Z(n8880) );
  MUX2_X2 U13450 ( .A(decode_regfile_intregs_2__1_), .B(
        decode_regfile_intregs_3__1_), .S(n10779), .Z(n8881) );
  MUX2_X2 U13451 ( .A(decode_regfile_intregs_0__1_), .B(
        decode_regfile_intregs_1__1_), .S(n10779), .Z(n8882) );
  MUX2_X2 U13452 ( .A(n8882), .B(n8881), .S(n10880), .Z(n8883) );
  MUX2_X2 U13453 ( .A(n8883), .B(n8880), .S(n10922), .Z(n8884) );
  MUX2_X2 U13454 ( .A(n8884), .B(n8877), .S(decode_rs2_3_), .Z(n8885) );
  MUX2_X2 U13455 ( .A(n8885), .B(n8870), .S(decode_rs2_4_), .Z(
        decode_regfile_N90) );
  MUX2_X2 U13456 ( .A(decode_regfile_intregs_30__2_), .B(
        decode_regfile_intregs_31__2_), .S(n10779), .Z(n8886) );
  MUX2_X2 U13457 ( .A(decode_regfile_intregs_28__2_), .B(
        decode_regfile_intregs_29__2_), .S(n10779), .Z(n8887) );
  MUX2_X2 U13458 ( .A(n8887), .B(n8886), .S(n10880), .Z(n8888) );
  MUX2_X2 U13459 ( .A(decode_regfile_intregs_26__2_), .B(
        decode_regfile_intregs_27__2_), .S(n10780), .Z(n8889) );
  MUX2_X2 U13460 ( .A(decode_regfile_intregs_24__2_), .B(
        decode_regfile_intregs_25__2_), .S(n10780), .Z(n8890) );
  MUX2_X2 U13461 ( .A(n8890), .B(n8889), .S(n10881), .Z(n8891) );
  MUX2_X2 U13462 ( .A(n8891), .B(n8888), .S(n10922), .Z(n8892) );
  MUX2_X2 U13463 ( .A(decode_regfile_intregs_22__2_), .B(
        decode_regfile_intregs_23__2_), .S(n10780), .Z(n8893) );
  MUX2_X2 U13464 ( .A(decode_regfile_intregs_20__2_), .B(
        decode_regfile_intregs_21__2_), .S(n10780), .Z(n8894) );
  MUX2_X2 U13465 ( .A(n8894), .B(n8893), .S(n10881), .Z(n8895) );
  MUX2_X2 U13466 ( .A(decode_regfile_intregs_18__2_), .B(
        decode_regfile_intregs_19__2_), .S(n10780), .Z(n8896) );
  MUX2_X2 U13467 ( .A(decode_regfile_intregs_16__2_), .B(
        decode_regfile_intregs_17__2_), .S(n10780), .Z(n8897) );
  MUX2_X2 U13468 ( .A(n8897), .B(n8896), .S(n10881), .Z(n8898) );
  MUX2_X2 U13469 ( .A(n8898), .B(n8895), .S(n10922), .Z(n8899) );
  MUX2_X2 U13470 ( .A(n8899), .B(n8892), .S(decode_rs2_3_), .Z(n8900) );
  MUX2_X2 U13471 ( .A(decode_regfile_intregs_14__2_), .B(
        decode_regfile_intregs_15__2_), .S(n10780), .Z(n8901) );
  MUX2_X2 U13472 ( .A(decode_regfile_intregs_12__2_), .B(
        decode_regfile_intregs_13__2_), .S(n10780), .Z(n8902) );
  MUX2_X2 U13473 ( .A(n8902), .B(n8901), .S(n10881), .Z(n8903) );
  MUX2_X2 U13474 ( .A(decode_regfile_intregs_10__2_), .B(
        decode_regfile_intregs_11__2_), .S(n10780), .Z(n8904) );
  MUX2_X2 U13475 ( .A(decode_regfile_intregs_8__2_), .B(
        decode_regfile_intregs_9__2_), .S(n10780), .Z(n8905) );
  MUX2_X2 U13476 ( .A(n8905), .B(n8904), .S(n10881), .Z(n8906) );
  MUX2_X2 U13477 ( .A(n8906), .B(n8903), .S(n10922), .Z(n8907) );
  MUX2_X2 U13478 ( .A(decode_regfile_intregs_6__2_), .B(
        decode_regfile_intregs_7__2_), .S(n10780), .Z(n8908) );
  MUX2_X2 U13479 ( .A(decode_regfile_intregs_4__2_), .B(
        decode_regfile_intregs_5__2_), .S(n10781), .Z(n8909) );
  MUX2_X2 U13480 ( .A(n8909), .B(n8908), .S(n10881), .Z(n8910) );
  MUX2_X2 U13481 ( .A(decode_regfile_intregs_2__2_), .B(
        decode_regfile_intregs_3__2_), .S(n10781), .Z(n8911) );
  MUX2_X2 U13482 ( .A(decode_regfile_intregs_0__2_), .B(
        decode_regfile_intregs_1__2_), .S(n10781), .Z(n8912) );
  MUX2_X2 U13483 ( .A(n8912), .B(n8911), .S(n10881), .Z(n8913) );
  MUX2_X2 U13484 ( .A(n8913), .B(n8910), .S(n10922), .Z(n8914) );
  MUX2_X2 U13485 ( .A(n8914), .B(n8907), .S(decode_rs2_3_), .Z(n8915) );
  MUX2_X2 U13486 ( .A(n8915), .B(n8900), .S(decode_rs2_4_), .Z(
        decode_regfile_N89) );
  MUX2_X2 U13487 ( .A(decode_regfile_intregs_30__3_), .B(
        decode_regfile_intregs_31__3_), .S(n10781), .Z(n8916) );
  MUX2_X2 U13488 ( .A(decode_regfile_intregs_28__3_), .B(
        decode_regfile_intregs_29__3_), .S(n10781), .Z(n8917) );
  MUX2_X2 U13489 ( .A(n8917), .B(n8916), .S(n10881), .Z(n8918) );
  MUX2_X2 U13490 ( .A(decode_regfile_intregs_26__3_), .B(
        decode_regfile_intregs_27__3_), .S(n10781), .Z(n8919) );
  MUX2_X2 U13491 ( .A(decode_regfile_intregs_24__3_), .B(
        decode_regfile_intregs_25__3_), .S(n10781), .Z(n8920) );
  MUX2_X2 U13492 ( .A(n8920), .B(n8919), .S(n10881), .Z(n8921) );
  MUX2_X2 U13493 ( .A(n8921), .B(n8918), .S(n10922), .Z(n8922) );
  MUX2_X2 U13494 ( .A(decode_regfile_intregs_22__3_), .B(
        decode_regfile_intregs_23__3_), .S(n10781), .Z(n8923) );
  MUX2_X2 U13495 ( .A(decode_regfile_intregs_20__3_), .B(
        decode_regfile_intregs_21__3_), .S(n10781), .Z(n8924) );
  MUX2_X2 U13496 ( .A(n8924), .B(n8923), .S(n10881), .Z(n8925) );
  MUX2_X2 U13497 ( .A(decode_regfile_intregs_18__3_), .B(
        decode_regfile_intregs_19__3_), .S(n10781), .Z(n8926) );
  MUX2_X2 U13498 ( .A(decode_regfile_intregs_16__3_), .B(
        decode_regfile_intregs_17__3_), .S(n10781), .Z(n8927) );
  MUX2_X2 U13499 ( .A(n8927), .B(n8926), .S(n10881), .Z(n8928) );
  MUX2_X2 U13500 ( .A(n8928), .B(n8925), .S(n10922), .Z(n8929) );
  MUX2_X2 U13501 ( .A(n8929), .B(n8922), .S(decode_rs2_3_), .Z(n8930) );
  MUX2_X2 U13502 ( .A(decode_regfile_intregs_14__3_), .B(
        decode_regfile_intregs_15__3_), .S(n10782), .Z(n8931) );
  MUX2_X2 U13503 ( .A(decode_regfile_intregs_12__3_), .B(
        decode_regfile_intregs_13__3_), .S(n10782), .Z(n8932) );
  MUX2_X2 U13504 ( .A(n8932), .B(n8931), .S(n10882), .Z(n8933) );
  MUX2_X2 U13505 ( .A(decode_regfile_intregs_10__3_), .B(
        decode_regfile_intregs_11__3_), .S(n10782), .Z(n8934) );
  MUX2_X2 U13506 ( .A(decode_regfile_intregs_8__3_), .B(
        decode_regfile_intregs_9__3_), .S(n10782), .Z(n8935) );
  MUX2_X2 U13507 ( .A(n8935), .B(n8934), .S(n10882), .Z(n8936) );
  MUX2_X2 U13508 ( .A(n8936), .B(n8933), .S(n10923), .Z(n8937) );
  MUX2_X2 U13509 ( .A(decode_regfile_intregs_6__3_), .B(
        decode_regfile_intregs_7__3_), .S(n10782), .Z(n8938) );
  MUX2_X2 U13510 ( .A(decode_regfile_intregs_4__3_), .B(
        decode_regfile_intregs_5__3_), .S(n10782), .Z(n8939) );
  MUX2_X2 U13511 ( .A(n8939), .B(n8938), .S(n10882), .Z(n8940) );
  MUX2_X2 U13512 ( .A(decode_regfile_intregs_2__3_), .B(
        decode_regfile_intregs_3__3_), .S(n10782), .Z(n8941) );
  MUX2_X2 U13513 ( .A(decode_regfile_intregs_0__3_), .B(
        decode_regfile_intregs_1__3_), .S(n10782), .Z(n8942) );
  MUX2_X2 U13514 ( .A(n8942), .B(n8941), .S(n10882), .Z(n8943) );
  MUX2_X2 U13515 ( .A(n8943), .B(n8940), .S(n10923), .Z(n8944) );
  MUX2_X2 U13516 ( .A(n8944), .B(n8937), .S(n10944), .Z(n8945) );
  MUX2_X2 U13517 ( .A(n8945), .B(n8930), .S(decode_rs2_4_), .Z(
        decode_regfile_N88) );
  MUX2_X2 U13518 ( .A(decode_regfile_intregs_30__4_), .B(
        decode_regfile_intregs_31__4_), .S(n10782), .Z(n8946) );
  MUX2_X2 U13519 ( .A(decode_regfile_intregs_28__4_), .B(
        decode_regfile_intregs_29__4_), .S(n10782), .Z(n8947) );
  MUX2_X2 U13520 ( .A(n8947), .B(n8946), .S(n10882), .Z(n8948) );
  MUX2_X2 U13521 ( .A(decode_regfile_intregs_26__4_), .B(
        decode_regfile_intregs_27__4_), .S(n10782), .Z(n8949) );
  MUX2_X2 U13522 ( .A(decode_regfile_intregs_24__4_), .B(
        decode_regfile_intregs_25__4_), .S(n10783), .Z(n8950) );
  MUX2_X2 U13523 ( .A(n8950), .B(n8949), .S(n10882), .Z(n8951) );
  MUX2_X2 U13524 ( .A(n8951), .B(n8948), .S(n10923), .Z(n8952) );
  MUX2_X2 U13525 ( .A(decode_regfile_intregs_22__4_), .B(
        decode_regfile_intregs_23__4_), .S(n10783), .Z(n8953) );
  MUX2_X2 U13526 ( .A(decode_regfile_intregs_20__4_), .B(
        decode_regfile_intregs_21__4_), .S(n10783), .Z(n8954) );
  MUX2_X2 U13527 ( .A(n8954), .B(n8953), .S(n10882), .Z(n8955) );
  MUX2_X2 U13528 ( .A(decode_regfile_intregs_18__4_), .B(
        decode_regfile_intregs_19__4_), .S(n10783), .Z(n8956) );
  MUX2_X2 U13529 ( .A(decode_regfile_intregs_16__4_), .B(
        decode_regfile_intregs_17__4_), .S(n10783), .Z(n8957) );
  MUX2_X2 U13530 ( .A(n8957), .B(n8956), .S(n10882), .Z(n8958) );
  MUX2_X2 U13531 ( .A(n8958), .B(n8955), .S(n10923), .Z(n8959) );
  MUX2_X2 U13532 ( .A(n8959), .B(n8952), .S(n10944), .Z(n8960) );
  MUX2_X2 U13533 ( .A(decode_regfile_intregs_14__4_), .B(
        decode_regfile_intregs_15__4_), .S(n10783), .Z(n8961) );
  MUX2_X2 U13534 ( .A(decode_regfile_intregs_12__4_), .B(
        decode_regfile_intregs_13__4_), .S(n10783), .Z(n8962) );
  MUX2_X2 U13535 ( .A(n8962), .B(n8961), .S(n10882), .Z(n8963) );
  MUX2_X2 U13536 ( .A(decode_regfile_intregs_10__4_), .B(
        decode_regfile_intregs_11__4_), .S(n10783), .Z(n8964) );
  MUX2_X2 U13537 ( .A(decode_regfile_intregs_8__4_), .B(
        decode_regfile_intregs_9__4_), .S(n10783), .Z(n8965) );
  MUX2_X2 U13538 ( .A(n8965), .B(n8964), .S(n10882), .Z(n8966) );
  MUX2_X2 U13539 ( .A(n8966), .B(n8963), .S(n10923), .Z(n8967) );
  MUX2_X2 U13540 ( .A(decode_regfile_intregs_6__4_), .B(
        decode_regfile_intregs_7__4_), .S(n10783), .Z(n8968) );
  MUX2_X2 U13541 ( .A(decode_regfile_intregs_4__4_), .B(
        decode_regfile_intregs_5__4_), .S(n10783), .Z(n8969) );
  MUX2_X2 U13542 ( .A(n8969), .B(n8968), .S(n10882), .Z(n8970) );
  MUX2_X2 U13543 ( .A(decode_regfile_intregs_2__4_), .B(
        decode_regfile_intregs_3__4_), .S(n10784), .Z(n8971) );
  MUX2_X2 U13544 ( .A(decode_regfile_intregs_0__4_), .B(
        decode_regfile_intregs_1__4_), .S(n10784), .Z(n8972) );
  MUX2_X2 U13545 ( .A(n8972), .B(n8971), .S(n10883), .Z(n8973) );
  MUX2_X2 U13546 ( .A(n8973), .B(n8970), .S(n10923), .Z(n8974) );
  MUX2_X2 U13547 ( .A(n8974), .B(n8967), .S(n10944), .Z(n8975) );
  MUX2_X2 U13548 ( .A(n8975), .B(n8960), .S(decode_rs2_4_), .Z(
        decode_regfile_N87) );
  MUX2_X2 U13549 ( .A(decode_regfile_intregs_30__5_), .B(
        decode_regfile_intregs_31__5_), .S(n10784), .Z(n8976) );
  MUX2_X2 U13550 ( .A(decode_regfile_intregs_28__5_), .B(
        decode_regfile_intregs_29__5_), .S(n10784), .Z(n8977) );
  MUX2_X2 U13551 ( .A(n8977), .B(n8976), .S(n10883), .Z(n8978) );
  MUX2_X2 U13552 ( .A(decode_regfile_intregs_26__5_), .B(
        decode_regfile_intregs_27__5_), .S(n10784), .Z(n8979) );
  MUX2_X2 U13553 ( .A(decode_regfile_intregs_24__5_), .B(
        decode_regfile_intregs_25__5_), .S(n10784), .Z(n8980) );
  MUX2_X2 U13554 ( .A(n8980), .B(n8979), .S(n10883), .Z(n8981) );
  MUX2_X2 U13555 ( .A(n8981), .B(n8978), .S(n10923), .Z(n8982) );
  MUX2_X2 U13556 ( .A(decode_regfile_intregs_22__5_), .B(
        decode_regfile_intregs_23__5_), .S(n10784), .Z(n8983) );
  MUX2_X2 U13557 ( .A(decode_regfile_intregs_20__5_), .B(
        decode_regfile_intregs_21__5_), .S(n10784), .Z(n8984) );
  MUX2_X2 U13558 ( .A(n8984), .B(n8983), .S(n10883), .Z(n8985) );
  MUX2_X2 U13559 ( .A(decode_regfile_intregs_18__5_), .B(
        decode_regfile_intregs_19__5_), .S(n10784), .Z(n8986) );
  MUX2_X2 U13560 ( .A(decode_regfile_intregs_16__5_), .B(
        decode_regfile_intregs_17__5_), .S(n10784), .Z(n8987) );
  MUX2_X2 U13561 ( .A(n8987), .B(n8986), .S(n10883), .Z(n8988) );
  MUX2_X2 U13562 ( .A(n8988), .B(n8985), .S(n10923), .Z(n8989) );
  MUX2_X2 U13563 ( .A(n8989), .B(n8982), .S(n10944), .Z(n8990) );
  MUX2_X2 U13564 ( .A(decode_regfile_intregs_14__5_), .B(
        decode_regfile_intregs_15__5_), .S(n10784), .Z(n8991) );
  MUX2_X2 U13565 ( .A(decode_regfile_intregs_12__5_), .B(
        decode_regfile_intregs_13__5_), .S(n10785), .Z(n8992) );
  MUX2_X2 U13566 ( .A(n8992), .B(n8991), .S(n10883), .Z(n8993) );
  MUX2_X2 U13567 ( .A(decode_regfile_intregs_10__5_), .B(
        decode_regfile_intregs_11__5_), .S(n10785), .Z(n8994) );
  MUX2_X2 U13568 ( .A(decode_regfile_intregs_8__5_), .B(
        decode_regfile_intregs_9__5_), .S(n10785), .Z(n8995) );
  MUX2_X2 U13569 ( .A(n8995), .B(n8994), .S(n10883), .Z(n8996) );
  MUX2_X2 U13570 ( .A(n8996), .B(n8993), .S(n10923), .Z(n8997) );
  MUX2_X2 U13571 ( .A(decode_regfile_intregs_6__5_), .B(
        decode_regfile_intregs_7__5_), .S(n10785), .Z(n8998) );
  MUX2_X2 U13572 ( .A(decode_regfile_intregs_4__5_), .B(
        decode_regfile_intregs_5__5_), .S(n10785), .Z(n8999) );
  MUX2_X2 U13573 ( .A(n8999), .B(n8998), .S(n10883), .Z(n9000) );
  MUX2_X2 U13574 ( .A(decode_regfile_intregs_2__5_), .B(
        decode_regfile_intregs_3__5_), .S(n10785), .Z(n9001) );
  MUX2_X2 U13575 ( .A(decode_regfile_intregs_0__5_), .B(
        decode_regfile_intregs_1__5_), .S(n10785), .Z(n9002) );
  MUX2_X2 U13576 ( .A(n9002), .B(n9001), .S(n10883), .Z(n9003) );
  MUX2_X2 U13577 ( .A(n9003), .B(n9000), .S(n10923), .Z(n9004) );
  MUX2_X2 U13578 ( .A(n9004), .B(n8997), .S(n10944), .Z(n9005) );
  MUX2_X2 U13579 ( .A(n9005), .B(n8990), .S(decode_rs2_4_), .Z(
        decode_regfile_N86) );
  MUX2_X2 U13580 ( .A(decode_regfile_intregs_30__6_), .B(
        decode_regfile_intregs_31__6_), .S(n10785), .Z(n9006) );
  MUX2_X2 U13581 ( .A(decode_regfile_intregs_28__6_), .B(
        decode_regfile_intregs_29__6_), .S(n10785), .Z(n9007) );
  MUX2_X2 U13582 ( .A(n9007), .B(n9006), .S(n10883), .Z(n9008) );
  MUX2_X2 U13583 ( .A(decode_regfile_intregs_26__6_), .B(
        decode_regfile_intregs_27__6_), .S(n10785), .Z(n9009) );
  MUX2_X2 U13584 ( .A(decode_regfile_intregs_24__6_), .B(
        decode_regfile_intregs_25__6_), .S(n10785), .Z(n9010) );
  MUX2_X2 U13585 ( .A(n9010), .B(n9009), .S(n10883), .Z(n9011) );
  MUX2_X2 U13586 ( .A(n9011), .B(n9008), .S(n10923), .Z(n9012) );
  MUX2_X2 U13587 ( .A(decode_regfile_intregs_22__6_), .B(
        decode_regfile_intregs_23__6_), .S(n10786), .Z(n9013) );
  MUX2_X2 U13588 ( .A(decode_regfile_intregs_20__6_), .B(
        decode_regfile_intregs_21__6_), .S(n10786), .Z(n9014) );
  MUX2_X2 U13589 ( .A(n9014), .B(n9013), .S(n10884), .Z(n9015) );
  MUX2_X2 U13590 ( .A(decode_regfile_intregs_18__6_), .B(
        decode_regfile_intregs_19__6_), .S(n10786), .Z(n9016) );
  MUX2_X2 U13591 ( .A(decode_regfile_intregs_16__6_), .B(
        decode_regfile_intregs_17__6_), .S(n10786), .Z(n9017) );
  MUX2_X2 U13592 ( .A(n9017), .B(n9016), .S(n10884), .Z(n9018) );
  MUX2_X2 U13593 ( .A(n9018), .B(n9015), .S(n10924), .Z(n9019) );
  MUX2_X2 U13594 ( .A(n9019), .B(n9012), .S(n10944), .Z(n9020) );
  MUX2_X2 U13595 ( .A(decode_regfile_intregs_14__6_), .B(
        decode_regfile_intregs_15__6_), .S(n10786), .Z(n9021) );
  MUX2_X2 U13596 ( .A(decode_regfile_intregs_12__6_), .B(
        decode_regfile_intregs_13__6_), .S(n10786), .Z(n9022) );
  MUX2_X2 U13597 ( .A(n9022), .B(n9021), .S(n10884), .Z(n9023) );
  MUX2_X2 U13598 ( .A(decode_regfile_intregs_10__6_), .B(
        decode_regfile_intregs_11__6_), .S(n10786), .Z(n9024) );
  MUX2_X2 U13599 ( .A(decode_regfile_intregs_8__6_), .B(
        decode_regfile_intregs_9__6_), .S(n10786), .Z(n9025) );
  MUX2_X2 U13600 ( .A(n9025), .B(n9024), .S(n10884), .Z(n9026) );
  MUX2_X2 U13601 ( .A(n9026), .B(n9023), .S(n10924), .Z(n9027) );
  MUX2_X2 U13602 ( .A(decode_regfile_intregs_6__6_), .B(
        decode_regfile_intregs_7__6_), .S(n10786), .Z(n9028) );
  MUX2_X2 U13603 ( .A(decode_regfile_intregs_4__6_), .B(
        decode_regfile_intregs_5__6_), .S(n10786), .Z(n9029) );
  MUX2_X2 U13604 ( .A(n9029), .B(n9028), .S(n10884), .Z(n9030) );
  MUX2_X2 U13605 ( .A(decode_regfile_intregs_2__6_), .B(
        decode_regfile_intregs_3__6_), .S(n10786), .Z(n9031) );
  MUX2_X2 U13606 ( .A(decode_regfile_intregs_0__6_), .B(
        decode_regfile_intregs_1__6_), .S(n10787), .Z(n9032) );
  MUX2_X2 U13607 ( .A(n9032), .B(n9031), .S(n10884), .Z(n9033) );
  MUX2_X2 U13608 ( .A(n9033), .B(n9030), .S(n10924), .Z(n9034) );
  MUX2_X2 U13609 ( .A(n9034), .B(n9027), .S(n10944), .Z(n9035) );
  MUX2_X2 U13610 ( .A(n9035), .B(n9020), .S(decode_rs2_4_), .Z(
        decode_regfile_N85) );
  MUX2_X2 U13611 ( .A(decode_regfile_intregs_30__7_), .B(
        decode_regfile_intregs_31__7_), .S(n10787), .Z(n9036) );
  MUX2_X2 U13612 ( .A(decode_regfile_intregs_28__7_), .B(
        decode_regfile_intregs_29__7_), .S(n10787), .Z(n9037) );
  MUX2_X2 U13613 ( .A(n9037), .B(n9036), .S(n10884), .Z(n9038) );
  MUX2_X2 U13614 ( .A(decode_regfile_intregs_26__7_), .B(
        decode_regfile_intregs_27__7_), .S(n10787), .Z(n9039) );
  MUX2_X2 U13615 ( .A(decode_regfile_intregs_24__7_), .B(
        decode_regfile_intregs_25__7_), .S(n10787), .Z(n9040) );
  MUX2_X2 U13616 ( .A(n9040), .B(n9039), .S(n10884), .Z(n9041) );
  MUX2_X2 U13617 ( .A(n9041), .B(n9038), .S(n10924), .Z(n9042) );
  MUX2_X2 U13618 ( .A(decode_regfile_intregs_22__7_), .B(
        decode_regfile_intregs_23__7_), .S(n10787), .Z(n9043) );
  MUX2_X2 U13619 ( .A(decode_regfile_intregs_20__7_), .B(
        decode_regfile_intregs_21__7_), .S(n10787), .Z(n9044) );
  MUX2_X2 U13620 ( .A(n9044), .B(n9043), .S(n10884), .Z(n9045) );
  MUX2_X2 U13621 ( .A(decode_regfile_intregs_18__7_), .B(
        decode_regfile_intregs_19__7_), .S(n10787), .Z(n9046) );
  MUX2_X2 U13622 ( .A(decode_regfile_intregs_16__7_), .B(
        decode_regfile_intregs_17__7_), .S(n10787), .Z(n9047) );
  MUX2_X2 U13623 ( .A(n9047), .B(n9046), .S(n10884), .Z(n9048) );
  MUX2_X2 U13624 ( .A(n9048), .B(n9045), .S(n10924), .Z(n9049) );
  MUX2_X2 U13625 ( .A(n9049), .B(n9042), .S(n10944), .Z(n9050) );
  MUX2_X2 U13626 ( .A(decode_regfile_intregs_14__7_), .B(
        decode_regfile_intregs_15__7_), .S(n10787), .Z(n9051) );
  MUX2_X2 U13627 ( .A(decode_regfile_intregs_12__7_), .B(
        decode_regfile_intregs_13__7_), .S(n10787), .Z(n9052) );
  MUX2_X2 U13628 ( .A(n9052), .B(n9051), .S(n10884), .Z(n9053) );
  MUX2_X2 U13629 ( .A(decode_regfile_intregs_10__7_), .B(
        decode_regfile_intregs_11__7_), .S(n10788), .Z(n9054) );
  MUX2_X2 U13630 ( .A(decode_regfile_intregs_8__7_), .B(
        decode_regfile_intregs_9__7_), .S(n10788), .Z(n9055) );
  MUX2_X2 U13631 ( .A(n9055), .B(n9054), .S(n10885), .Z(n9056) );
  MUX2_X2 U13632 ( .A(n9056), .B(n9053), .S(n10924), .Z(n9057) );
  MUX2_X2 U13633 ( .A(decode_regfile_intregs_6__7_), .B(
        decode_regfile_intregs_7__7_), .S(n10788), .Z(n9058) );
  MUX2_X2 U13634 ( .A(decode_regfile_intregs_4__7_), .B(
        decode_regfile_intregs_5__7_), .S(n10788), .Z(n9059) );
  MUX2_X2 U13635 ( .A(n9059), .B(n9058), .S(n10885), .Z(n9060) );
  MUX2_X2 U13636 ( .A(decode_regfile_intregs_2__7_), .B(
        decode_regfile_intregs_3__7_), .S(n10788), .Z(n9061) );
  MUX2_X2 U13637 ( .A(decode_regfile_intregs_0__7_), .B(
        decode_regfile_intregs_1__7_), .S(n10788), .Z(n9062) );
  MUX2_X2 U13638 ( .A(n9062), .B(n9061), .S(n10885), .Z(n9063) );
  MUX2_X2 U13639 ( .A(n9063), .B(n9060), .S(n10924), .Z(n9064) );
  MUX2_X2 U13640 ( .A(n9064), .B(n9057), .S(n10944), .Z(n9065) );
  MUX2_X2 U13641 ( .A(n9065), .B(n9050), .S(decode_rs2_4_), .Z(
        decode_regfile_N84) );
  MUX2_X2 U13642 ( .A(decode_regfile_intregs_30__8_), .B(
        decode_regfile_intregs_31__8_), .S(n10788), .Z(n9066) );
  MUX2_X2 U13643 ( .A(decode_regfile_intregs_28__8_), .B(
        decode_regfile_intregs_29__8_), .S(n10788), .Z(n9067) );
  MUX2_X2 U13644 ( .A(n9067), .B(n9066), .S(n10885), .Z(n9068) );
  MUX2_X2 U13645 ( .A(decode_regfile_intregs_26__8_), .B(
        decode_regfile_intregs_27__8_), .S(n10788), .Z(n9069) );
  MUX2_X2 U13646 ( .A(decode_regfile_intregs_24__8_), .B(
        decode_regfile_intregs_25__8_), .S(n10788), .Z(n9070) );
  MUX2_X2 U13647 ( .A(n9070), .B(n9069), .S(n10885), .Z(n9071) );
  MUX2_X2 U13648 ( .A(n9071), .B(n9068), .S(n10924), .Z(n9072) );
  MUX2_X2 U13649 ( .A(decode_regfile_intregs_22__8_), .B(
        decode_regfile_intregs_23__8_), .S(n10788), .Z(n9073) );
  MUX2_X2 U13650 ( .A(decode_regfile_intregs_20__8_), .B(
        decode_regfile_intregs_21__8_), .S(n10789), .Z(n9074) );
  MUX2_X2 U13651 ( .A(n9074), .B(n9073), .S(n10885), .Z(n9075) );
  MUX2_X2 U13652 ( .A(decode_regfile_intregs_18__8_), .B(
        decode_regfile_intregs_19__8_), .S(n10789), .Z(n9076) );
  MUX2_X2 U13653 ( .A(decode_regfile_intregs_16__8_), .B(
        decode_regfile_intregs_17__8_), .S(n10789), .Z(n9077) );
  MUX2_X2 U13654 ( .A(n9077), .B(n9076), .S(n10885), .Z(n9078) );
  MUX2_X2 U13655 ( .A(n9078), .B(n9075), .S(n10924), .Z(n9079) );
  MUX2_X2 U13656 ( .A(n9079), .B(n9072), .S(n10944), .Z(n9080) );
  MUX2_X2 U13657 ( .A(decode_regfile_intregs_14__8_), .B(
        decode_regfile_intregs_15__8_), .S(n10789), .Z(n9081) );
  MUX2_X2 U13658 ( .A(decode_regfile_intregs_12__8_), .B(
        decode_regfile_intregs_13__8_), .S(n10789), .Z(n9082) );
  MUX2_X2 U13659 ( .A(n9082), .B(n9081), .S(n10885), .Z(n9083) );
  MUX2_X2 U13660 ( .A(decode_regfile_intregs_10__8_), .B(
        decode_regfile_intregs_11__8_), .S(n10789), .Z(n9084) );
  MUX2_X2 U13661 ( .A(decode_regfile_intregs_8__8_), .B(
        decode_regfile_intregs_9__8_), .S(n10789), .Z(n9085) );
  MUX2_X2 U13662 ( .A(n9085), .B(n9084), .S(n10885), .Z(n9086) );
  MUX2_X2 U13663 ( .A(n9086), .B(n9083), .S(n10924), .Z(n9087) );
  MUX2_X2 U13664 ( .A(decode_regfile_intregs_6__8_), .B(
        decode_regfile_intregs_7__8_), .S(n10789), .Z(n9088) );
  MUX2_X2 U13665 ( .A(decode_regfile_intregs_4__8_), .B(
        decode_regfile_intregs_5__8_), .S(n10789), .Z(n9089) );
  MUX2_X2 U13666 ( .A(n9089), .B(n9088), .S(n10885), .Z(n9090) );
  MUX2_X2 U13667 ( .A(decode_regfile_intregs_2__8_), .B(
        decode_regfile_intregs_3__8_), .S(n10789), .Z(n9091) );
  MUX2_X2 U13668 ( .A(decode_regfile_intregs_0__8_), .B(
        decode_regfile_intregs_1__8_), .S(n10789), .Z(n9092) );
  MUX2_X2 U13669 ( .A(n9092), .B(n9091), .S(n10885), .Z(n9093) );
  MUX2_X2 U13670 ( .A(n9093), .B(n9090), .S(n10924), .Z(n9094) );
  MUX2_X2 U13671 ( .A(n9094), .B(n9087), .S(n10944), .Z(n9095) );
  MUX2_X2 U13672 ( .A(n9095), .B(n9080), .S(decode_rs2_4_), .Z(
        decode_regfile_N83) );
  MUX2_X2 U13673 ( .A(decode_regfile_intregs_30__9_), .B(
        decode_regfile_intregs_31__9_), .S(n10790), .Z(n9096) );
  MUX2_X2 U13674 ( .A(decode_regfile_intregs_28__9_), .B(
        decode_regfile_intregs_29__9_), .S(n10790), .Z(n9097) );
  MUX2_X2 U13675 ( .A(n9097), .B(n9096), .S(n10886), .Z(n9098) );
  MUX2_X2 U13676 ( .A(decode_regfile_intregs_26__9_), .B(
        decode_regfile_intregs_27__9_), .S(n10790), .Z(n9099) );
  MUX2_X2 U13677 ( .A(decode_regfile_intregs_24__9_), .B(
        decode_regfile_intregs_25__9_), .S(n10790), .Z(n9100) );
  MUX2_X2 U13678 ( .A(n9100), .B(n9099), .S(n10886), .Z(n9101) );
  MUX2_X2 U13679 ( .A(n9101), .B(n9098), .S(n10925), .Z(n9102) );
  MUX2_X2 U13680 ( .A(decode_regfile_intregs_22__9_), .B(
        decode_regfile_intregs_23__9_), .S(n10790), .Z(n9103) );
  MUX2_X2 U13681 ( .A(decode_regfile_intregs_20__9_), .B(
        decode_regfile_intregs_21__9_), .S(n10790), .Z(n9104) );
  MUX2_X2 U13682 ( .A(n9104), .B(n9103), .S(n10886), .Z(n9105) );
  MUX2_X2 U13683 ( .A(decode_regfile_intregs_18__9_), .B(
        decode_regfile_intregs_19__9_), .S(n10790), .Z(n9106) );
  MUX2_X2 U13684 ( .A(decode_regfile_intregs_16__9_), .B(
        decode_regfile_intregs_17__9_), .S(n10790), .Z(n9107) );
  MUX2_X2 U13685 ( .A(n9107), .B(n9106), .S(n10886), .Z(n9108) );
  MUX2_X2 U13686 ( .A(n9108), .B(n9105), .S(n10925), .Z(n9109) );
  MUX2_X2 U13687 ( .A(n9109), .B(n9102), .S(n10945), .Z(n9110) );
  MUX2_X2 U13688 ( .A(decode_regfile_intregs_14__9_), .B(
        decode_regfile_intregs_15__9_), .S(n10790), .Z(n9111) );
  MUX2_X2 U13689 ( .A(decode_regfile_intregs_12__9_), .B(
        decode_regfile_intregs_13__9_), .S(n10790), .Z(n9112) );
  MUX2_X2 U13690 ( .A(n9112), .B(n9111), .S(n10886), .Z(n9113) );
  MUX2_X2 U13691 ( .A(decode_regfile_intregs_10__9_), .B(
        decode_regfile_intregs_11__9_), .S(n10790), .Z(n9114) );
  MUX2_X2 U13692 ( .A(decode_regfile_intregs_8__9_), .B(
        decode_regfile_intregs_9__9_), .S(n10791), .Z(n9115) );
  MUX2_X2 U13693 ( .A(n9115), .B(n9114), .S(n10886), .Z(n9116) );
  MUX2_X2 U13694 ( .A(n9116), .B(n9113), .S(n10925), .Z(n9117) );
  MUX2_X2 U13695 ( .A(decode_regfile_intregs_6__9_), .B(
        decode_regfile_intregs_7__9_), .S(n10791), .Z(n9118) );
  MUX2_X2 U13696 ( .A(decode_regfile_intregs_4__9_), .B(
        decode_regfile_intregs_5__9_), .S(n10791), .Z(n9119) );
  MUX2_X2 U13697 ( .A(n9119), .B(n9118), .S(n10886), .Z(n9120) );
  MUX2_X2 U13698 ( .A(decode_regfile_intregs_2__9_), .B(
        decode_regfile_intregs_3__9_), .S(n10791), .Z(n9121) );
  MUX2_X2 U13699 ( .A(decode_regfile_intregs_0__9_), .B(
        decode_regfile_intregs_1__9_), .S(n10791), .Z(n9122) );
  MUX2_X2 U13700 ( .A(n9122), .B(n9121), .S(n10886), .Z(n9123) );
  MUX2_X2 U13701 ( .A(n9123), .B(n9120), .S(n10925), .Z(n9124) );
  MUX2_X2 U13702 ( .A(n9124), .B(n9117), .S(n10945), .Z(n9125) );
  MUX2_X2 U13703 ( .A(n9125), .B(n9110), .S(n10956), .Z(decode_regfile_N82) );
  MUX2_X2 U13704 ( .A(decode_regfile_intregs_30__10_), .B(
        decode_regfile_intregs_31__10_), .S(n10791), .Z(n9126) );
  MUX2_X2 U13705 ( .A(decode_regfile_intregs_28__10_), .B(
        decode_regfile_intregs_29__10_), .S(n10791), .Z(n9127) );
  MUX2_X2 U13706 ( .A(n9127), .B(n9126), .S(n10886), .Z(n9128) );
  MUX2_X2 U13707 ( .A(decode_regfile_intregs_26__10_), .B(
        decode_regfile_intregs_27__10_), .S(n10791), .Z(n9129) );
  MUX2_X2 U13708 ( .A(decode_regfile_intregs_24__10_), .B(
        decode_regfile_intregs_25__10_), .S(n10791), .Z(n9130) );
  MUX2_X2 U13709 ( .A(n9130), .B(n9129), .S(n10886), .Z(n9131) );
  MUX2_X2 U13710 ( .A(n9131), .B(n9128), .S(n10925), .Z(n9132) );
  MUX2_X2 U13711 ( .A(decode_regfile_intregs_22__10_), .B(
        decode_regfile_intregs_23__10_), .S(n10791), .Z(n9133) );
  MUX2_X2 U13712 ( .A(decode_regfile_intregs_20__10_), .B(
        decode_regfile_intregs_21__10_), .S(n10791), .Z(n9134) );
  MUX2_X2 U13713 ( .A(n9134), .B(n9133), .S(n10886), .Z(n9135) );
  MUX2_X2 U13714 ( .A(decode_regfile_intregs_18__10_), .B(
        decode_regfile_intregs_19__10_), .S(n10792), .Z(n9136) );
  MUX2_X2 U13715 ( .A(decode_regfile_intregs_16__10_), .B(
        decode_regfile_intregs_17__10_), .S(n10792), .Z(n9137) );
  MUX2_X2 U13716 ( .A(n9137), .B(n9136), .S(n10887), .Z(n9138) );
  MUX2_X2 U13717 ( .A(n9138), .B(n9135), .S(n10925), .Z(n9139) );
  MUX2_X2 U13718 ( .A(n9139), .B(n9132), .S(n10945), .Z(n9140) );
  MUX2_X2 U13719 ( .A(decode_regfile_intregs_14__10_), .B(
        decode_regfile_intregs_15__10_), .S(n10792), .Z(n9141) );
  MUX2_X2 U13720 ( .A(decode_regfile_intregs_12__10_), .B(
        decode_regfile_intregs_13__10_), .S(n10792), .Z(n9142) );
  MUX2_X2 U13721 ( .A(n9142), .B(n9141), .S(n10887), .Z(n9143) );
  MUX2_X2 U13722 ( .A(decode_regfile_intregs_10__10_), .B(
        decode_regfile_intregs_11__10_), .S(n10792), .Z(n9144) );
  MUX2_X2 U13723 ( .A(decode_regfile_intregs_8__10_), .B(
        decode_regfile_intregs_9__10_), .S(n10792), .Z(n9145) );
  MUX2_X2 U13724 ( .A(n9145), .B(n9144), .S(n10887), .Z(n9146) );
  MUX2_X2 U13725 ( .A(n9146), .B(n9143), .S(n10925), .Z(n9147) );
  MUX2_X2 U13726 ( .A(decode_regfile_intregs_6__10_), .B(
        decode_regfile_intregs_7__10_), .S(n10792), .Z(n9148) );
  MUX2_X2 U13727 ( .A(decode_regfile_intregs_4__10_), .B(
        decode_regfile_intregs_5__10_), .S(n10792), .Z(n9149) );
  MUX2_X2 U13728 ( .A(n9149), .B(n9148), .S(n10887), .Z(n9150) );
  MUX2_X2 U13729 ( .A(decode_regfile_intregs_2__10_), .B(
        decode_regfile_intregs_3__10_), .S(n10792), .Z(n9151) );
  MUX2_X2 U13730 ( .A(decode_regfile_intregs_0__10_), .B(
        decode_regfile_intregs_1__10_), .S(n10792), .Z(n9152) );
  MUX2_X2 U13731 ( .A(n9152), .B(n9151), .S(n10887), .Z(n9153) );
  MUX2_X2 U13732 ( .A(n9153), .B(n9150), .S(n10925), .Z(n9154) );
  MUX2_X2 U13733 ( .A(n9154), .B(n9147), .S(n10945), .Z(n9155) );
  MUX2_X2 U13734 ( .A(n9155), .B(n9140), .S(n10956), .Z(decode_regfile_N81) );
  MUX2_X2 U13735 ( .A(decode_regfile_intregs_30__11_), .B(
        decode_regfile_intregs_31__11_), .S(n10792), .Z(n9156) );
  MUX2_X2 U13736 ( .A(decode_regfile_intregs_28__11_), .B(
        decode_regfile_intregs_29__11_), .S(n10793), .Z(n9157) );
  MUX2_X2 U13737 ( .A(n9157), .B(n9156), .S(n10887), .Z(n9158) );
  MUX2_X2 U13738 ( .A(decode_regfile_intregs_26__11_), .B(
        decode_regfile_intregs_27__11_), .S(n10793), .Z(n9159) );
  MUX2_X2 U13739 ( .A(decode_regfile_intregs_24__11_), .B(
        decode_regfile_intregs_25__11_), .S(n10793), .Z(n9160) );
  MUX2_X2 U13740 ( .A(n9160), .B(n9159), .S(n10887), .Z(n9161) );
  MUX2_X2 U13741 ( .A(n9161), .B(n9158), .S(n10925), .Z(n9162) );
  MUX2_X2 U13742 ( .A(decode_regfile_intregs_22__11_), .B(
        decode_regfile_intregs_23__11_), .S(n10793), .Z(n9163) );
  MUX2_X2 U13743 ( .A(decode_regfile_intregs_20__11_), .B(
        decode_regfile_intregs_21__11_), .S(n10793), .Z(n9164) );
  MUX2_X2 U13744 ( .A(n9164), .B(n9163), .S(n10887), .Z(n9165) );
  MUX2_X2 U13745 ( .A(decode_regfile_intregs_18__11_), .B(
        decode_regfile_intregs_19__11_), .S(n10793), .Z(n9166) );
  MUX2_X2 U13746 ( .A(decode_regfile_intregs_16__11_), .B(
        decode_regfile_intregs_17__11_), .S(n10793), .Z(n9167) );
  MUX2_X2 U13747 ( .A(n9167), .B(n9166), .S(n10887), .Z(n9168) );
  MUX2_X2 U13748 ( .A(n9168), .B(n9165), .S(n10925), .Z(n9169) );
  MUX2_X2 U13749 ( .A(n9169), .B(n9162), .S(n10945), .Z(n9170) );
  MUX2_X2 U13750 ( .A(decode_regfile_intregs_14__11_), .B(
        decode_regfile_intregs_15__11_), .S(n10793), .Z(n9171) );
  MUX2_X2 U13751 ( .A(decode_regfile_intregs_12__11_), .B(
        decode_regfile_intregs_13__11_), .S(n10793), .Z(n9172) );
  MUX2_X2 U13752 ( .A(n9172), .B(n9171), .S(n10887), .Z(n9173) );
  MUX2_X2 U13753 ( .A(decode_regfile_intregs_10__11_), .B(
        decode_regfile_intregs_11__11_), .S(n10793), .Z(n9174) );
  MUX2_X2 U13754 ( .A(decode_regfile_intregs_8__11_), .B(
        decode_regfile_intregs_9__11_), .S(n10793), .Z(n9175) );
  MUX2_X2 U13755 ( .A(n9175), .B(n9174), .S(n10887), .Z(n9176) );
  MUX2_X2 U13756 ( .A(n9176), .B(n9173), .S(n10925), .Z(n9177) );
  MUX2_X2 U13757 ( .A(decode_regfile_intregs_6__11_), .B(
        decode_regfile_intregs_7__11_), .S(n10794), .Z(n9178) );
  MUX2_X2 U13758 ( .A(decode_regfile_intregs_4__11_), .B(
        decode_regfile_intregs_5__11_), .S(n10794), .Z(n9179) );
  MUX2_X2 U13759 ( .A(n9179), .B(n9178), .S(n10888), .Z(n9180) );
  MUX2_X2 U13760 ( .A(decode_regfile_intregs_2__11_), .B(
        decode_regfile_intregs_3__11_), .S(n10794), .Z(n9181) );
  MUX2_X2 U13761 ( .A(decode_regfile_intregs_0__11_), .B(
        decode_regfile_intregs_1__11_), .S(n10794), .Z(n9182) );
  MUX2_X2 U13762 ( .A(n9182), .B(n9181), .S(n10888), .Z(n9183) );
  MUX2_X2 U13763 ( .A(n9183), .B(n9180), .S(n10926), .Z(n9184) );
  MUX2_X2 U13764 ( .A(n9184), .B(n9177), .S(n10945), .Z(n9185) );
  MUX2_X2 U13765 ( .A(n9185), .B(n9170), .S(n10956), .Z(decode_regfile_N80) );
  MUX2_X2 U13766 ( .A(decode_regfile_intregs_30__12_), .B(
        decode_regfile_intregs_31__12_), .S(n10794), .Z(n9186) );
  MUX2_X2 U13767 ( .A(decode_regfile_intregs_28__12_), .B(
        decode_regfile_intregs_29__12_), .S(n10794), .Z(n9187) );
  MUX2_X2 U13768 ( .A(n9187), .B(n9186), .S(n10888), .Z(n9188) );
  MUX2_X2 U13769 ( .A(decode_regfile_intregs_26__12_), .B(
        decode_regfile_intregs_27__12_), .S(n10794), .Z(n9189) );
  MUX2_X2 U13770 ( .A(decode_regfile_intregs_24__12_), .B(
        decode_regfile_intregs_25__12_), .S(n10794), .Z(n9190) );
  MUX2_X2 U13771 ( .A(n9190), .B(n9189), .S(n10888), .Z(n9191) );
  MUX2_X2 U13772 ( .A(n9191), .B(n9188), .S(n10926), .Z(n9192) );
  MUX2_X2 U13773 ( .A(decode_regfile_intregs_22__12_), .B(
        decode_regfile_intregs_23__12_), .S(n10794), .Z(n9193) );
  MUX2_X2 U13774 ( .A(decode_regfile_intregs_20__12_), .B(
        decode_regfile_intregs_21__12_), .S(n10794), .Z(n9194) );
  MUX2_X2 U13775 ( .A(n9194), .B(n9193), .S(n10888), .Z(n9195) );
  MUX2_X2 U13776 ( .A(decode_regfile_intregs_18__12_), .B(
        decode_regfile_intregs_19__12_), .S(n10794), .Z(n9196) );
  MUX2_X2 U13777 ( .A(decode_regfile_intregs_16__12_), .B(
        decode_regfile_intregs_17__12_), .S(n10795), .Z(n9197) );
  MUX2_X2 U13778 ( .A(n9197), .B(n9196), .S(n10888), .Z(n9198) );
  MUX2_X2 U13779 ( .A(n9198), .B(n9195), .S(n10926), .Z(n9199) );
  MUX2_X2 U13780 ( .A(n9199), .B(n9192), .S(n10945), .Z(n9200) );
  MUX2_X2 U13781 ( .A(decode_regfile_intregs_14__12_), .B(
        decode_regfile_intregs_15__12_), .S(n10795), .Z(n9201) );
  MUX2_X2 U13782 ( .A(decode_regfile_intregs_12__12_), .B(
        decode_regfile_intregs_13__12_), .S(n10795), .Z(n9202) );
  MUX2_X2 U13783 ( .A(n9202), .B(n9201), .S(n10888), .Z(n9203) );
  MUX2_X2 U13784 ( .A(decode_regfile_intregs_10__12_), .B(
        decode_regfile_intregs_11__12_), .S(n10795), .Z(n9204) );
  MUX2_X2 U13785 ( .A(decode_regfile_intregs_8__12_), .B(
        decode_regfile_intregs_9__12_), .S(n10795), .Z(n9205) );
  MUX2_X2 U13786 ( .A(n9205), .B(n9204), .S(n10888), .Z(n9206) );
  MUX2_X2 U13787 ( .A(n9206), .B(n9203), .S(n10926), .Z(n9207) );
  MUX2_X2 U13788 ( .A(decode_regfile_intregs_6__12_), .B(
        decode_regfile_intregs_7__12_), .S(n10795), .Z(n9208) );
  MUX2_X2 U13789 ( .A(decode_regfile_intregs_4__12_), .B(
        decode_regfile_intregs_5__12_), .S(n10795), .Z(n9209) );
  MUX2_X2 U13790 ( .A(n9209), .B(n9208), .S(n10888), .Z(n9210) );
  MUX2_X2 U13791 ( .A(decode_regfile_intregs_2__12_), .B(
        decode_regfile_intregs_3__12_), .S(n10795), .Z(n9211) );
  MUX2_X2 U13792 ( .A(decode_regfile_intregs_0__12_), .B(
        decode_regfile_intregs_1__12_), .S(n10795), .Z(n9212) );
  MUX2_X2 U13793 ( .A(n9212), .B(n9211), .S(n10888), .Z(n9213) );
  MUX2_X2 U13794 ( .A(n9213), .B(n9210), .S(n10926), .Z(n9214) );
  MUX2_X2 U13795 ( .A(n9214), .B(n9207), .S(n10945), .Z(n9215) );
  MUX2_X2 U13796 ( .A(n9215), .B(n9200), .S(n10956), .Z(decode_regfile_N79) );
  MUX2_X2 U13797 ( .A(decode_regfile_intregs_30__13_), .B(
        decode_regfile_intregs_31__13_), .S(n10795), .Z(n9216) );
  MUX2_X2 U13798 ( .A(decode_regfile_intregs_28__13_), .B(
        decode_regfile_intregs_29__13_), .S(n10795), .Z(n9217) );
  MUX2_X2 U13799 ( .A(n9217), .B(n9216), .S(n10888), .Z(n9218) );
  MUX2_X2 U13800 ( .A(decode_regfile_intregs_26__13_), .B(
        decode_regfile_intregs_27__13_), .S(n10796), .Z(n9219) );
  MUX2_X2 U13801 ( .A(decode_regfile_intregs_24__13_), .B(
        decode_regfile_intregs_25__13_), .S(n10796), .Z(n9220) );
  MUX2_X2 U13802 ( .A(n9220), .B(n9219), .S(n10889), .Z(n9221) );
  MUX2_X2 U13803 ( .A(n9221), .B(n9218), .S(n10926), .Z(n9222) );
  MUX2_X2 U13804 ( .A(decode_regfile_intregs_22__13_), .B(
        decode_regfile_intregs_23__13_), .S(n10796), .Z(n9223) );
  MUX2_X2 U13805 ( .A(decode_regfile_intregs_20__13_), .B(
        decode_regfile_intregs_21__13_), .S(n10796), .Z(n9224) );
  MUX2_X2 U13806 ( .A(n9224), .B(n9223), .S(n10889), .Z(n9225) );
  MUX2_X2 U13807 ( .A(decode_regfile_intregs_18__13_), .B(
        decode_regfile_intregs_19__13_), .S(n10796), .Z(n9226) );
  MUX2_X2 U13808 ( .A(decode_regfile_intregs_16__13_), .B(
        decode_regfile_intregs_17__13_), .S(n10796), .Z(n9227) );
  MUX2_X2 U13809 ( .A(n9227), .B(n9226), .S(n10889), .Z(n9228) );
  MUX2_X2 U13810 ( .A(n9228), .B(n9225), .S(n10926), .Z(n9229) );
  MUX2_X2 U13811 ( .A(n9229), .B(n9222), .S(n10945), .Z(n9230) );
  MUX2_X2 U13812 ( .A(decode_regfile_intregs_14__13_), .B(
        decode_regfile_intregs_15__13_), .S(n10796), .Z(n9231) );
  MUX2_X2 U13813 ( .A(decode_regfile_intregs_12__13_), .B(
        decode_regfile_intregs_13__13_), .S(n10796), .Z(n9232) );
  MUX2_X2 U13814 ( .A(n9232), .B(n9231), .S(n10889), .Z(n9233) );
  MUX2_X2 U13815 ( .A(decode_regfile_intregs_10__13_), .B(
        decode_regfile_intregs_11__13_), .S(n10796), .Z(n9234) );
  MUX2_X2 U13816 ( .A(decode_regfile_intregs_8__13_), .B(
        decode_regfile_intregs_9__13_), .S(n10796), .Z(n9235) );
  MUX2_X2 U13817 ( .A(n9235), .B(n9234), .S(n10889), .Z(n9236) );
  MUX2_X2 U13818 ( .A(n9236), .B(n9233), .S(n10926), .Z(n9237) );
  MUX2_X2 U13819 ( .A(decode_regfile_intregs_6__13_), .B(
        decode_regfile_intregs_7__13_), .S(n10796), .Z(n9238) );
  MUX2_X2 U13820 ( .A(decode_regfile_intregs_4__13_), .B(
        decode_regfile_intregs_5__13_), .S(n10797), .Z(n9239) );
  MUX2_X2 U13821 ( .A(n9239), .B(n9238), .S(n10889), .Z(n9240) );
  MUX2_X2 U13822 ( .A(decode_regfile_intregs_2__13_), .B(
        decode_regfile_intregs_3__13_), .S(n10797), .Z(n9241) );
  MUX2_X2 U13823 ( .A(decode_regfile_intregs_0__13_), .B(
        decode_regfile_intregs_1__13_), .S(n10797), .Z(n9242) );
  MUX2_X2 U13824 ( .A(n9242), .B(n9241), .S(n10889), .Z(n9243) );
  MUX2_X2 U13825 ( .A(n9243), .B(n9240), .S(n10926), .Z(n9244) );
  MUX2_X2 U13826 ( .A(n9244), .B(n9237), .S(n10945), .Z(n9245) );
  MUX2_X2 U13827 ( .A(n9245), .B(n9230), .S(n10956), .Z(decode_regfile_N78) );
  MUX2_X2 U13828 ( .A(decode_regfile_intregs_30__14_), .B(
        decode_regfile_intregs_31__14_), .S(n10797), .Z(n9246) );
  MUX2_X2 U13829 ( .A(decode_regfile_intregs_28__14_), .B(
        decode_regfile_intregs_29__14_), .S(n10797), .Z(n9247) );
  MUX2_X2 U13830 ( .A(n9247), .B(n9246), .S(n10889), .Z(n9248) );
  MUX2_X2 U13831 ( .A(decode_regfile_intregs_26__14_), .B(
        decode_regfile_intregs_27__14_), .S(n10797), .Z(n9249) );
  MUX2_X2 U13832 ( .A(decode_regfile_intregs_24__14_), .B(
        decode_regfile_intregs_25__14_), .S(n10797), .Z(n9250) );
  MUX2_X2 U13833 ( .A(n9250), .B(n9249), .S(n10889), .Z(n9251) );
  MUX2_X2 U13834 ( .A(n9251), .B(n9248), .S(n10926), .Z(n9252) );
  MUX2_X2 U13835 ( .A(decode_regfile_intregs_22__14_), .B(
        decode_regfile_intregs_23__14_), .S(n10797), .Z(n9253) );
  MUX2_X2 U13836 ( .A(decode_regfile_intregs_20__14_), .B(
        decode_regfile_intregs_21__14_), .S(n10797), .Z(n9254) );
  MUX2_X2 U13837 ( .A(n9254), .B(n9253), .S(n10889), .Z(n9255) );
  MUX2_X2 U13838 ( .A(decode_regfile_intregs_18__14_), .B(
        decode_regfile_intregs_19__14_), .S(n10797), .Z(n9256) );
  MUX2_X2 U13839 ( .A(decode_regfile_intregs_16__14_), .B(
        decode_regfile_intregs_17__14_), .S(n10797), .Z(n9257) );
  MUX2_X2 U13840 ( .A(n9257), .B(n9256), .S(n10889), .Z(n9258) );
  MUX2_X2 U13841 ( .A(n9258), .B(n9255), .S(n10926), .Z(n9259) );
  MUX2_X2 U13842 ( .A(n9259), .B(n9252), .S(n10945), .Z(n9260) );
  MUX2_X2 U13843 ( .A(decode_regfile_intregs_14__14_), .B(
        decode_regfile_intregs_15__14_), .S(n10798), .Z(n9261) );
  MUX2_X2 U13844 ( .A(decode_regfile_intregs_12__14_), .B(
        decode_regfile_intregs_13__14_), .S(n10798), .Z(n9262) );
  MUX2_X2 U13845 ( .A(n9262), .B(n9261), .S(n10890), .Z(n9263) );
  MUX2_X2 U13846 ( .A(decode_regfile_intregs_10__14_), .B(
        decode_regfile_intregs_11__14_), .S(n10798), .Z(n9264) );
  MUX2_X2 U13847 ( .A(decode_regfile_intregs_8__14_), .B(
        decode_regfile_intregs_9__14_), .S(n10798), .Z(n9265) );
  MUX2_X2 U13848 ( .A(n9265), .B(n9264), .S(n10890), .Z(n9266) );
  MUX2_X2 U13849 ( .A(n9266), .B(n9263), .S(n10927), .Z(n9267) );
  MUX2_X2 U13850 ( .A(decode_regfile_intregs_6__14_), .B(
        decode_regfile_intregs_7__14_), .S(n10798), .Z(n9268) );
  MUX2_X2 U13851 ( .A(decode_regfile_intregs_4__14_), .B(
        decode_regfile_intregs_5__14_), .S(n10798), .Z(n9269) );
  MUX2_X2 U13852 ( .A(n9269), .B(n9268), .S(n10890), .Z(n9270) );
  MUX2_X2 U13853 ( .A(decode_regfile_intregs_2__14_), .B(
        decode_regfile_intregs_3__14_), .S(n10798), .Z(n9271) );
  MUX2_X2 U13854 ( .A(decode_regfile_intregs_0__14_), .B(
        decode_regfile_intregs_1__14_), .S(n10798), .Z(n9272) );
  MUX2_X2 U13855 ( .A(n9272), .B(n9271), .S(n10890), .Z(n9273) );
  MUX2_X2 U13856 ( .A(n9273), .B(n9270), .S(n10927), .Z(n9274) );
  MUX2_X2 U13857 ( .A(n9274), .B(n9267), .S(n10946), .Z(n9275) );
  MUX2_X2 U13858 ( .A(n9275), .B(n9260), .S(n10956), .Z(decode_regfile_N77) );
  MUX2_X2 U13859 ( .A(decode_regfile_intregs_30__15_), .B(
        decode_regfile_intregs_31__15_), .S(n10798), .Z(n9276) );
  MUX2_X2 U13860 ( .A(decode_regfile_intregs_28__15_), .B(
        decode_regfile_intregs_29__15_), .S(n10798), .Z(n9277) );
  MUX2_X2 U13861 ( .A(n9277), .B(n9276), .S(n10890), .Z(n9278) );
  MUX2_X2 U13862 ( .A(decode_regfile_intregs_26__15_), .B(
        decode_regfile_intregs_27__15_), .S(n10798), .Z(n9279) );
  MUX2_X2 U13863 ( .A(decode_regfile_intregs_24__15_), .B(
        decode_regfile_intregs_25__15_), .S(n10799), .Z(n9280) );
  MUX2_X2 U13864 ( .A(n9280), .B(n9279), .S(n10890), .Z(n9281) );
  MUX2_X2 U13865 ( .A(n9281), .B(n9278), .S(n10927), .Z(n9282) );
  MUX2_X2 U13866 ( .A(decode_regfile_intregs_22__15_), .B(
        decode_regfile_intregs_23__15_), .S(n10799), .Z(n9283) );
  MUX2_X2 U13867 ( .A(decode_regfile_intregs_20__15_), .B(
        decode_regfile_intregs_21__15_), .S(n10799), .Z(n9284) );
  MUX2_X2 U13868 ( .A(n9284), .B(n9283), .S(n10890), .Z(n9285) );
  MUX2_X2 U13869 ( .A(decode_regfile_intregs_18__15_), .B(
        decode_regfile_intregs_19__15_), .S(n10799), .Z(n9286) );
  MUX2_X2 U13870 ( .A(decode_regfile_intregs_16__15_), .B(
        decode_regfile_intregs_17__15_), .S(n10799), .Z(n9287) );
  MUX2_X2 U13871 ( .A(n9287), .B(n9286), .S(n10890), .Z(n9288) );
  MUX2_X2 U13872 ( .A(n9288), .B(n9285), .S(n10927), .Z(n9289) );
  MUX2_X2 U13873 ( .A(n9289), .B(n9282), .S(n10946), .Z(n9290) );
  MUX2_X2 U13874 ( .A(decode_regfile_intregs_14__15_), .B(
        decode_regfile_intregs_15__15_), .S(n10799), .Z(n9291) );
  MUX2_X2 U13875 ( .A(decode_regfile_intregs_12__15_), .B(
        decode_regfile_intregs_13__15_), .S(n10799), .Z(n9292) );
  MUX2_X2 U13876 ( .A(n9292), .B(n9291), .S(n10890), .Z(n9293) );
  MUX2_X2 U13877 ( .A(decode_regfile_intregs_10__15_), .B(
        decode_regfile_intregs_11__15_), .S(n10799), .Z(n9294) );
  MUX2_X2 U13878 ( .A(decode_regfile_intregs_8__15_), .B(
        decode_regfile_intregs_9__15_), .S(n10799), .Z(n9295) );
  MUX2_X2 U13879 ( .A(n9295), .B(n9294), .S(n10890), .Z(n9296) );
  MUX2_X2 U13880 ( .A(n9296), .B(n9293), .S(n10927), .Z(n9297) );
  MUX2_X2 U13881 ( .A(decode_regfile_intregs_6__15_), .B(
        decode_regfile_intregs_7__15_), .S(n10799), .Z(n9298) );
  MUX2_X2 U13882 ( .A(decode_regfile_intregs_4__15_), .B(
        decode_regfile_intregs_5__15_), .S(n10799), .Z(n9299) );
  MUX2_X2 U13883 ( .A(n9299), .B(n9298), .S(n10890), .Z(n9300) );
  MUX2_X2 U13884 ( .A(decode_regfile_intregs_2__15_), .B(
        decode_regfile_intregs_3__15_), .S(n10800), .Z(n9301) );
  MUX2_X2 U13885 ( .A(decode_regfile_intregs_0__15_), .B(
        decode_regfile_intregs_1__15_), .S(n10800), .Z(n9302) );
  MUX2_X2 U13886 ( .A(n9302), .B(n9301), .S(n10891), .Z(n9303) );
  MUX2_X2 U13887 ( .A(n9303), .B(n9300), .S(n10927), .Z(n9304) );
  MUX2_X2 U13888 ( .A(n9304), .B(n9297), .S(n10946), .Z(n9305) );
  MUX2_X2 U13889 ( .A(n9305), .B(n9290), .S(n10956), .Z(decode_regfile_N76) );
  MUX2_X2 U13890 ( .A(decode_regfile_intregs_30__16_), .B(
        decode_regfile_intregs_31__16_), .S(n10800), .Z(n9306) );
  MUX2_X2 U13891 ( .A(decode_regfile_intregs_28__16_), .B(
        decode_regfile_intregs_29__16_), .S(n10800), .Z(n9307) );
  MUX2_X2 U13892 ( .A(n9307), .B(n9306), .S(n10891), .Z(n9308) );
  MUX2_X2 U13893 ( .A(decode_regfile_intregs_26__16_), .B(
        decode_regfile_intregs_27__16_), .S(n10800), .Z(n9309) );
  MUX2_X2 U13894 ( .A(decode_regfile_intregs_24__16_), .B(
        decode_regfile_intregs_25__16_), .S(n10800), .Z(n9310) );
  MUX2_X2 U13895 ( .A(n9310), .B(n9309), .S(n10891), .Z(n9311) );
  MUX2_X2 U13896 ( .A(n9311), .B(n9308), .S(n10927), .Z(n9312) );
  MUX2_X2 U13897 ( .A(decode_regfile_intregs_22__16_), .B(
        decode_regfile_intregs_23__16_), .S(n10800), .Z(n9313) );
  MUX2_X2 U13898 ( .A(decode_regfile_intregs_20__16_), .B(
        decode_regfile_intregs_21__16_), .S(n10800), .Z(n9314) );
  MUX2_X2 U13899 ( .A(n9314), .B(n9313), .S(n10891), .Z(n9315) );
  MUX2_X2 U13900 ( .A(decode_regfile_intregs_18__16_), .B(
        decode_regfile_intregs_19__16_), .S(n10800), .Z(n9316) );
  MUX2_X2 U13901 ( .A(decode_regfile_intregs_16__16_), .B(
        decode_regfile_intregs_17__16_), .S(n10800), .Z(n9317) );
  MUX2_X2 U13902 ( .A(n9317), .B(n9316), .S(n10891), .Z(n9318) );
  MUX2_X2 U13903 ( .A(n9318), .B(n9315), .S(n10927), .Z(n9319) );
  MUX2_X2 U13904 ( .A(n9319), .B(n9312), .S(n10946), .Z(n9320) );
  MUX2_X2 U13905 ( .A(decode_regfile_intregs_14__16_), .B(
        decode_regfile_intregs_15__16_), .S(n10800), .Z(n9321) );
  MUX2_X2 U13906 ( .A(decode_regfile_intregs_12__16_), .B(
        decode_regfile_intregs_13__16_), .S(n10801), .Z(n9322) );
  MUX2_X2 U13907 ( .A(n9322), .B(n9321), .S(n10891), .Z(n9323) );
  MUX2_X2 U13908 ( .A(decode_regfile_intregs_10__16_), .B(
        decode_regfile_intregs_11__16_), .S(n10801), .Z(n9324) );
  MUX2_X2 U13909 ( .A(decode_regfile_intregs_8__16_), .B(
        decode_regfile_intregs_9__16_), .S(n10801), .Z(n9325) );
  MUX2_X2 U13910 ( .A(n9325), .B(n9324), .S(n10891), .Z(n9326) );
  MUX2_X2 U13911 ( .A(n9326), .B(n9323), .S(n10927), .Z(n9327) );
  MUX2_X2 U13912 ( .A(decode_regfile_intregs_6__16_), .B(
        decode_regfile_intregs_7__16_), .S(n10801), .Z(n9328) );
  MUX2_X2 U13913 ( .A(decode_regfile_intregs_4__16_), .B(
        decode_regfile_intregs_5__16_), .S(n10801), .Z(n9329) );
  MUX2_X2 U13914 ( .A(n9329), .B(n9328), .S(n10891), .Z(n9330) );
  MUX2_X2 U13915 ( .A(decode_regfile_intregs_2__16_), .B(
        decode_regfile_intregs_3__16_), .S(n10801), .Z(n9331) );
  MUX2_X2 U13916 ( .A(decode_regfile_intregs_0__16_), .B(
        decode_regfile_intregs_1__16_), .S(n10801), .Z(n9332) );
  MUX2_X2 U13917 ( .A(n9332), .B(n9331), .S(n10891), .Z(n9333) );
  MUX2_X2 U13918 ( .A(n9333), .B(n9330), .S(n10927), .Z(n9334) );
  MUX2_X2 U13919 ( .A(n9334), .B(n9327), .S(n10946), .Z(n9335) );
  MUX2_X2 U13920 ( .A(n9335), .B(n9320), .S(n10956), .Z(decode_regfile_N75) );
  MUX2_X2 U13921 ( .A(decode_regfile_intregs_30__17_), .B(
        decode_regfile_intregs_31__17_), .S(n10801), .Z(n9336) );
  MUX2_X2 U13922 ( .A(decode_regfile_intregs_28__17_), .B(
        decode_regfile_intregs_29__17_), .S(n10801), .Z(n9337) );
  MUX2_X2 U13923 ( .A(n9337), .B(n9336), .S(n10891), .Z(n9338) );
  MUX2_X2 U13924 ( .A(decode_regfile_intregs_26__17_), .B(
        decode_regfile_intregs_27__17_), .S(n10801), .Z(n9339) );
  MUX2_X2 U13925 ( .A(decode_regfile_intregs_24__17_), .B(
        decode_regfile_intregs_25__17_), .S(n10801), .Z(n9340) );
  MUX2_X2 U13926 ( .A(n9340), .B(n9339), .S(n10891), .Z(n9341) );
  MUX2_X2 U13927 ( .A(n9341), .B(n9338), .S(n10927), .Z(n9342) );
  MUX2_X2 U13928 ( .A(decode_regfile_intregs_22__17_), .B(
        decode_regfile_intregs_23__17_), .S(n10802), .Z(n9343) );
  MUX2_X2 U13929 ( .A(decode_regfile_intregs_20__17_), .B(
        decode_regfile_intregs_21__17_), .S(n10802), .Z(n9344) );
  MUX2_X2 U13930 ( .A(n9344), .B(n9343), .S(n10892), .Z(n9345) );
  MUX2_X2 U13931 ( .A(decode_regfile_intregs_18__17_), .B(
        decode_regfile_intregs_19__17_), .S(n10802), .Z(n9346) );
  MUX2_X2 U13932 ( .A(decode_regfile_intregs_16__17_), .B(
        decode_regfile_intregs_17__17_), .S(n10802), .Z(n9347) );
  MUX2_X2 U13933 ( .A(n9347), .B(n9346), .S(n10892), .Z(n9348) );
  MUX2_X2 U13934 ( .A(n9348), .B(n9345), .S(n10928), .Z(n9349) );
  MUX2_X2 U13935 ( .A(n9349), .B(n9342), .S(n10946), .Z(n9350) );
  MUX2_X2 U13936 ( .A(decode_regfile_intregs_14__17_), .B(
        decode_regfile_intregs_15__17_), .S(n10802), .Z(n9351) );
  MUX2_X2 U13937 ( .A(decode_regfile_intregs_12__17_), .B(
        decode_regfile_intregs_13__17_), .S(n10802), .Z(n9352) );
  MUX2_X2 U13938 ( .A(n9352), .B(n9351), .S(n10892), .Z(n9353) );
  MUX2_X2 U13939 ( .A(decode_regfile_intregs_10__17_), .B(
        decode_regfile_intregs_11__17_), .S(n10802), .Z(n9354) );
  MUX2_X2 U13940 ( .A(decode_regfile_intregs_8__17_), .B(
        decode_regfile_intregs_9__17_), .S(n10802), .Z(n9355) );
  MUX2_X2 U13941 ( .A(n9355), .B(n9354), .S(n10892), .Z(n9356) );
  MUX2_X2 U13942 ( .A(n9356), .B(n9353), .S(n10928), .Z(n9357) );
  MUX2_X2 U13943 ( .A(decode_regfile_intregs_6__17_), .B(
        decode_regfile_intregs_7__17_), .S(n10802), .Z(n9358) );
  MUX2_X2 U13944 ( .A(decode_regfile_intregs_4__17_), .B(
        decode_regfile_intregs_5__17_), .S(n10802), .Z(n9359) );
  MUX2_X2 U13945 ( .A(n9359), .B(n9358), .S(n10892), .Z(n9360) );
  MUX2_X2 U13946 ( .A(decode_regfile_intregs_2__17_), .B(
        decode_regfile_intregs_3__17_), .S(n10802), .Z(n9361) );
  MUX2_X2 U13947 ( .A(decode_regfile_intregs_0__17_), .B(
        decode_regfile_intregs_1__17_), .S(n10803), .Z(n9362) );
  MUX2_X2 U13948 ( .A(n9362), .B(n9361), .S(n10892), .Z(n9363) );
  MUX2_X2 U13949 ( .A(n9363), .B(n9360), .S(n10928), .Z(n9364) );
  MUX2_X2 U13950 ( .A(n9364), .B(n9357), .S(n10946), .Z(n9365) );
  MUX2_X2 U13951 ( .A(n9365), .B(n9350), .S(n10956), .Z(decode_regfile_N74) );
  MUX2_X2 U13952 ( .A(decode_regfile_intregs_30__18_), .B(
        decode_regfile_intregs_31__18_), .S(n10803), .Z(n9366) );
  MUX2_X2 U13953 ( .A(decode_regfile_intregs_28__18_), .B(
        decode_regfile_intregs_29__18_), .S(n10803), .Z(n9367) );
  MUX2_X2 U13954 ( .A(n9367), .B(n9366), .S(n10892), .Z(n9368) );
  MUX2_X2 U13955 ( .A(decode_regfile_intregs_26__18_), .B(
        decode_regfile_intregs_27__18_), .S(n10803), .Z(n9369) );
  MUX2_X2 U13956 ( .A(decode_regfile_intregs_24__18_), .B(
        decode_regfile_intregs_25__18_), .S(n10803), .Z(n9370) );
  MUX2_X2 U13957 ( .A(n9370), .B(n9369), .S(n10892), .Z(n9371) );
  MUX2_X2 U13958 ( .A(n9371), .B(n9368), .S(n10928), .Z(n9372) );
  MUX2_X2 U13959 ( .A(decode_regfile_intregs_22__18_), .B(
        decode_regfile_intregs_23__18_), .S(n10803), .Z(n9373) );
  MUX2_X2 U13960 ( .A(decode_regfile_intregs_20__18_), .B(
        decode_regfile_intregs_21__18_), .S(n10803), .Z(n9374) );
  MUX2_X2 U13961 ( .A(n9374), .B(n9373), .S(n10892), .Z(n9375) );
  MUX2_X2 U13962 ( .A(decode_regfile_intregs_18__18_), .B(
        decode_regfile_intregs_19__18_), .S(n10803), .Z(n9376) );
  MUX2_X2 U13963 ( .A(decode_regfile_intregs_16__18_), .B(
        decode_regfile_intregs_17__18_), .S(n10803), .Z(n9377) );
  MUX2_X2 U13964 ( .A(n9377), .B(n9376), .S(n10892), .Z(n9378) );
  MUX2_X2 U13965 ( .A(n9378), .B(n9375), .S(n10928), .Z(n9379) );
  MUX2_X2 U13966 ( .A(n9379), .B(n9372), .S(n10946), .Z(n9380) );
  MUX2_X2 U13967 ( .A(decode_regfile_intregs_14__18_), .B(
        decode_regfile_intregs_15__18_), .S(n10803), .Z(n9381) );
  MUX2_X2 U13968 ( .A(decode_regfile_intregs_12__18_), .B(
        decode_regfile_intregs_13__18_), .S(n10803), .Z(n9382) );
  MUX2_X2 U13969 ( .A(n9382), .B(n9381), .S(n10892), .Z(n9383) );
  MUX2_X2 U13970 ( .A(decode_regfile_intregs_10__18_), .B(
        decode_regfile_intregs_11__18_), .S(n10804), .Z(n9384) );
  MUX2_X2 U13971 ( .A(decode_regfile_intregs_8__18_), .B(
        decode_regfile_intregs_9__18_), .S(n10804), .Z(n9385) );
  MUX2_X2 U13972 ( .A(n9385), .B(n9384), .S(n10893), .Z(n9386) );
  MUX2_X2 U13973 ( .A(n9386), .B(n9383), .S(n10928), .Z(n9387) );
  MUX2_X2 U13974 ( .A(decode_regfile_intregs_6__18_), .B(
        decode_regfile_intregs_7__18_), .S(n10804), .Z(n9388) );
  MUX2_X2 U13975 ( .A(decode_regfile_intregs_4__18_), .B(
        decode_regfile_intregs_5__18_), .S(n10804), .Z(n9389) );
  MUX2_X2 U13976 ( .A(n9389), .B(n9388), .S(n10893), .Z(n9390) );
  MUX2_X2 U13977 ( .A(decode_regfile_intregs_2__18_), .B(
        decode_regfile_intregs_3__18_), .S(n10804), .Z(n9391) );
  MUX2_X2 U13978 ( .A(decode_regfile_intregs_0__18_), .B(
        decode_regfile_intregs_1__18_), .S(n10804), .Z(n9392) );
  MUX2_X2 U13979 ( .A(n9392), .B(n9391), .S(n10893), .Z(n9393) );
  MUX2_X2 U13980 ( .A(n9393), .B(n9390), .S(n10928), .Z(n9394) );
  MUX2_X2 U13981 ( .A(n9394), .B(n9387), .S(n10946), .Z(n9395) );
  MUX2_X2 U13982 ( .A(n9395), .B(n9380), .S(n10956), .Z(decode_regfile_N73) );
  MUX2_X2 U13983 ( .A(decode_regfile_intregs_30__19_), .B(
        decode_regfile_intregs_31__19_), .S(n10804), .Z(n9396) );
  MUX2_X2 U13984 ( .A(decode_regfile_intregs_28__19_), .B(
        decode_regfile_intregs_29__19_), .S(n10804), .Z(n9397) );
  MUX2_X2 U13985 ( .A(n9397), .B(n9396), .S(n10893), .Z(n9398) );
  MUX2_X2 U13986 ( .A(decode_regfile_intregs_26__19_), .B(
        decode_regfile_intregs_27__19_), .S(n10804), .Z(n9399) );
  MUX2_X2 U13987 ( .A(decode_regfile_intregs_24__19_), .B(
        decode_regfile_intregs_25__19_), .S(n10804), .Z(n9400) );
  MUX2_X2 U13988 ( .A(n9400), .B(n9399), .S(n10893), .Z(n9401) );
  MUX2_X2 U13989 ( .A(n9401), .B(n9398), .S(n10928), .Z(n9402) );
  MUX2_X2 U13990 ( .A(decode_regfile_intregs_22__19_), .B(
        decode_regfile_intregs_23__19_), .S(n10804), .Z(n9403) );
  MUX2_X2 U13991 ( .A(decode_regfile_intregs_20__19_), .B(
        decode_regfile_intregs_21__19_), .S(n10805), .Z(n9404) );
  MUX2_X2 U13992 ( .A(n9404), .B(n9403), .S(n10893), .Z(n9405) );
  MUX2_X2 U13993 ( .A(decode_regfile_intregs_18__19_), .B(
        decode_regfile_intregs_19__19_), .S(n10805), .Z(n9406) );
  MUX2_X2 U13994 ( .A(decode_regfile_intregs_16__19_), .B(
        decode_regfile_intregs_17__19_), .S(n10805), .Z(n9407) );
  MUX2_X2 U13995 ( .A(n9407), .B(n9406), .S(n10893), .Z(n9408) );
  MUX2_X2 U13996 ( .A(n9408), .B(n9405), .S(n10928), .Z(n9409) );
  MUX2_X2 U13997 ( .A(n9409), .B(n9402), .S(n10946), .Z(n9410) );
  MUX2_X2 U13998 ( .A(decode_regfile_intregs_14__19_), .B(
        decode_regfile_intregs_15__19_), .S(n10805), .Z(n9411) );
  MUX2_X2 U13999 ( .A(decode_regfile_intregs_12__19_), .B(
        decode_regfile_intregs_13__19_), .S(n10805), .Z(n9412) );
  MUX2_X2 U14000 ( .A(n9412), .B(n9411), .S(n10893), .Z(n9413) );
  MUX2_X2 U14001 ( .A(decode_regfile_intregs_10__19_), .B(
        decode_regfile_intregs_11__19_), .S(n10805), .Z(n9414) );
  MUX2_X2 U14002 ( .A(decode_regfile_intregs_8__19_), .B(
        decode_regfile_intregs_9__19_), .S(n10805), .Z(n9415) );
  MUX2_X2 U14003 ( .A(n9415), .B(n9414), .S(n10893), .Z(n9416) );
  MUX2_X2 U14004 ( .A(n9416), .B(n9413), .S(n10928), .Z(n9417) );
  MUX2_X2 U14005 ( .A(decode_regfile_intregs_6__19_), .B(
        decode_regfile_intregs_7__19_), .S(n10805), .Z(n9418) );
  MUX2_X2 U14006 ( .A(decode_regfile_intregs_4__19_), .B(
        decode_regfile_intregs_5__19_), .S(n10805), .Z(n9419) );
  MUX2_X2 U14007 ( .A(n9419), .B(n9418), .S(n10893), .Z(n9420) );
  MUX2_X2 U14008 ( .A(decode_regfile_intregs_2__19_), .B(
        decode_regfile_intregs_3__19_), .S(n10805), .Z(n9421) );
  MUX2_X2 U14009 ( .A(decode_regfile_intregs_0__19_), .B(
        decode_regfile_intregs_1__19_), .S(n10805), .Z(n9422) );
  MUX2_X2 U14010 ( .A(n9422), .B(n9421), .S(n10893), .Z(n9423) );
  MUX2_X2 U14011 ( .A(n9423), .B(n9420), .S(n10928), .Z(n9424) );
  MUX2_X2 U14012 ( .A(n9424), .B(n9417), .S(n10946), .Z(n9425) );
  MUX2_X2 U14013 ( .A(n9425), .B(n9410), .S(n10956), .Z(decode_regfile_N72) );
  MUX2_X2 U14014 ( .A(decode_regfile_intregs_30__20_), .B(
        decode_regfile_intregs_31__20_), .S(n10806), .Z(n9426) );
  MUX2_X2 U14015 ( .A(decode_regfile_intregs_28__20_), .B(
        decode_regfile_intregs_29__20_), .S(n10806), .Z(n9427) );
  MUX2_X2 U14016 ( .A(n9427), .B(n9426), .S(n10894), .Z(n9428) );
  MUX2_X2 U14017 ( .A(decode_regfile_intregs_26__20_), .B(
        decode_regfile_intregs_27__20_), .S(n10806), .Z(n9429) );
  MUX2_X2 U14018 ( .A(decode_regfile_intregs_24__20_), .B(
        decode_regfile_intregs_25__20_), .S(n10806), .Z(n9430) );
  MUX2_X2 U14019 ( .A(n9430), .B(n9429), .S(n10894), .Z(n9431) );
  MUX2_X2 U14020 ( .A(n9431), .B(n9428), .S(n10929), .Z(n9432) );
  MUX2_X2 U14021 ( .A(decode_regfile_intregs_22__20_), .B(
        decode_regfile_intregs_23__20_), .S(n10806), .Z(n9433) );
  MUX2_X2 U14022 ( .A(decode_regfile_intregs_20__20_), .B(
        decode_regfile_intregs_21__20_), .S(n10806), .Z(n9434) );
  MUX2_X2 U14023 ( .A(n9434), .B(n9433), .S(n10894), .Z(n9435) );
  MUX2_X2 U14024 ( .A(decode_regfile_intregs_18__20_), .B(
        decode_regfile_intregs_19__20_), .S(n10806), .Z(n9436) );
  MUX2_X2 U14025 ( .A(decode_regfile_intregs_16__20_), .B(
        decode_regfile_intregs_17__20_), .S(n10806), .Z(n9437) );
  MUX2_X2 U14026 ( .A(n9437), .B(n9436), .S(n10894), .Z(n9438) );
  MUX2_X2 U14027 ( .A(n9438), .B(n9435), .S(n10929), .Z(n9439) );
  MUX2_X2 U14028 ( .A(n9439), .B(n9432), .S(n10947), .Z(n9440) );
  MUX2_X2 U14029 ( .A(decode_regfile_intregs_14__20_), .B(
        decode_regfile_intregs_15__20_), .S(n10806), .Z(n9441) );
  MUX2_X2 U14030 ( .A(decode_regfile_intregs_12__20_), .B(
        decode_regfile_intregs_13__20_), .S(n10806), .Z(n9442) );
  MUX2_X2 U14031 ( .A(n9442), .B(n9441), .S(n10894), .Z(n9443) );
  MUX2_X2 U14032 ( .A(decode_regfile_intregs_10__20_), .B(
        decode_regfile_intregs_11__20_), .S(n10806), .Z(n9444) );
  MUX2_X2 U14033 ( .A(decode_regfile_intregs_8__20_), .B(
        decode_regfile_intregs_9__20_), .S(n10807), .Z(n9445) );
  MUX2_X2 U14034 ( .A(n9445), .B(n9444), .S(n10894), .Z(n9446) );
  MUX2_X2 U14035 ( .A(n9446), .B(n9443), .S(n10929), .Z(n9447) );
  MUX2_X2 U14036 ( .A(decode_regfile_intregs_6__20_), .B(
        decode_regfile_intregs_7__20_), .S(n10807), .Z(n9448) );
  MUX2_X2 U14037 ( .A(decode_regfile_intregs_4__20_), .B(
        decode_regfile_intregs_5__20_), .S(n10807), .Z(n9449) );
  MUX2_X2 U14038 ( .A(n9449), .B(n9448), .S(n10894), .Z(n9450) );
  MUX2_X2 U14039 ( .A(decode_regfile_intregs_2__20_), .B(
        decode_regfile_intregs_3__20_), .S(n10807), .Z(n9451) );
  MUX2_X2 U14040 ( .A(decode_regfile_intregs_0__20_), .B(
        decode_regfile_intregs_1__20_), .S(n10807), .Z(n9452) );
  MUX2_X2 U14041 ( .A(n9452), .B(n9451), .S(n10894), .Z(n9453) );
  MUX2_X2 U14042 ( .A(n9453), .B(n9450), .S(n10929), .Z(n9454) );
  MUX2_X2 U14043 ( .A(n9454), .B(n9447), .S(n10947), .Z(n9455) );
  MUX2_X2 U14044 ( .A(n9455), .B(n9440), .S(n10957), .Z(decode_regfile_N71) );
  MUX2_X2 U14045 ( .A(decode_regfile_intregs_30__21_), .B(
        decode_regfile_intregs_31__21_), .S(n10807), .Z(n9456) );
  MUX2_X2 U14046 ( .A(decode_regfile_intregs_28__21_), .B(
        decode_regfile_intregs_29__21_), .S(n10807), .Z(n9457) );
  MUX2_X2 U14047 ( .A(n9457), .B(n9456), .S(n10894), .Z(n9458) );
  MUX2_X2 U14048 ( .A(decode_regfile_intregs_26__21_), .B(
        decode_regfile_intregs_27__21_), .S(n10807), .Z(n9459) );
  MUX2_X2 U14049 ( .A(decode_regfile_intregs_24__21_), .B(
        decode_regfile_intregs_25__21_), .S(n10807), .Z(n9460) );
  MUX2_X2 U14050 ( .A(n9460), .B(n9459), .S(n10894), .Z(n9461) );
  MUX2_X2 U14051 ( .A(n9461), .B(n9458), .S(n10929), .Z(n9462) );
  MUX2_X2 U14052 ( .A(decode_regfile_intregs_22__21_), .B(
        decode_regfile_intregs_23__21_), .S(n10807), .Z(n9463) );
  MUX2_X2 U14053 ( .A(decode_regfile_intregs_20__21_), .B(
        decode_regfile_intregs_21__21_), .S(n10807), .Z(n9464) );
  MUX2_X2 U14054 ( .A(n9464), .B(n9463), .S(n10894), .Z(n9465) );
  MUX2_X2 U14055 ( .A(decode_regfile_intregs_18__21_), .B(
        decode_regfile_intregs_19__21_), .S(n10808), .Z(n9466) );
  MUX2_X2 U14056 ( .A(decode_regfile_intregs_16__21_), .B(
        decode_regfile_intregs_17__21_), .S(n10808), .Z(n9467) );
  MUX2_X2 U14057 ( .A(n9467), .B(n9466), .S(n10895), .Z(n9468) );
  MUX2_X2 U14058 ( .A(n9468), .B(n9465), .S(n10929), .Z(n9469) );
  MUX2_X2 U14059 ( .A(n9469), .B(n9462), .S(n10947), .Z(n9470) );
  MUX2_X2 U14060 ( .A(decode_regfile_intregs_14__21_), .B(
        decode_regfile_intregs_15__21_), .S(n10808), .Z(n9471) );
  MUX2_X2 U14061 ( .A(decode_regfile_intregs_12__21_), .B(
        decode_regfile_intregs_13__21_), .S(n10808), .Z(n9472) );
  MUX2_X2 U14062 ( .A(n9472), .B(n9471), .S(n10895), .Z(n9473) );
  MUX2_X2 U14063 ( .A(decode_regfile_intregs_10__21_), .B(
        decode_regfile_intregs_11__21_), .S(n10808), .Z(n9474) );
  MUX2_X2 U14064 ( .A(decode_regfile_intregs_8__21_), .B(
        decode_regfile_intregs_9__21_), .S(n10808), .Z(n9475) );
  MUX2_X2 U14065 ( .A(n9475), .B(n9474), .S(n10895), .Z(n9476) );
  MUX2_X2 U14066 ( .A(n9476), .B(n9473), .S(n10929), .Z(n9477) );
  MUX2_X2 U14067 ( .A(decode_regfile_intregs_6__21_), .B(
        decode_regfile_intregs_7__21_), .S(n10808), .Z(n9478) );
  MUX2_X2 U14068 ( .A(decode_regfile_intregs_4__21_), .B(
        decode_regfile_intregs_5__21_), .S(n10808), .Z(n9479) );
  MUX2_X2 U14069 ( .A(n9479), .B(n9478), .S(n10895), .Z(n9480) );
  MUX2_X2 U14070 ( .A(decode_regfile_intregs_2__21_), .B(
        decode_regfile_intregs_3__21_), .S(n10808), .Z(n9481) );
  MUX2_X2 U14071 ( .A(decode_regfile_intregs_0__21_), .B(
        decode_regfile_intregs_1__21_), .S(n10808), .Z(n9482) );
  MUX2_X2 U14072 ( .A(n9482), .B(n9481), .S(n10895), .Z(n9483) );
  MUX2_X2 U14073 ( .A(n9483), .B(n9480), .S(n10929), .Z(n9484) );
  MUX2_X2 U14074 ( .A(n9484), .B(n9477), .S(n10947), .Z(n9485) );
  MUX2_X2 U14075 ( .A(n9485), .B(n9470), .S(n10957), .Z(decode_regfile_N70) );
  MUX2_X2 U14076 ( .A(decode_regfile_intregs_30__22_), .B(
        decode_regfile_intregs_31__22_), .S(n10808), .Z(n9486) );
  MUX2_X2 U14077 ( .A(decode_regfile_intregs_28__22_), .B(
        decode_regfile_intregs_29__22_), .S(n10809), .Z(n9487) );
  MUX2_X2 U14078 ( .A(n9487), .B(n9486), .S(n10895), .Z(n9488) );
  MUX2_X2 U14079 ( .A(decode_regfile_intregs_26__22_), .B(
        decode_regfile_intregs_27__22_), .S(n10809), .Z(n9489) );
  MUX2_X2 U14080 ( .A(decode_regfile_intregs_24__22_), .B(
        decode_regfile_intregs_25__22_), .S(n10809), .Z(n9490) );
  MUX2_X2 U14081 ( .A(n9490), .B(n9489), .S(n10895), .Z(n9491) );
  MUX2_X2 U14082 ( .A(n9491), .B(n9488), .S(n10929), .Z(n9492) );
  MUX2_X2 U14083 ( .A(decode_regfile_intregs_22__22_), .B(
        decode_regfile_intregs_23__22_), .S(n10809), .Z(n9493) );
  MUX2_X2 U14084 ( .A(decode_regfile_intregs_20__22_), .B(
        decode_regfile_intregs_21__22_), .S(n10809), .Z(n9494) );
  MUX2_X2 U14085 ( .A(n9494), .B(n9493), .S(n10895), .Z(n9495) );
  MUX2_X2 U14086 ( .A(decode_regfile_intregs_18__22_), .B(
        decode_regfile_intregs_19__22_), .S(n10809), .Z(n9496) );
  MUX2_X2 U14087 ( .A(decode_regfile_intregs_16__22_), .B(
        decode_regfile_intregs_17__22_), .S(n10809), .Z(n9497) );
  MUX2_X2 U14088 ( .A(n9497), .B(n9496), .S(n10895), .Z(n9498) );
  MUX2_X2 U14089 ( .A(n9498), .B(n9495), .S(n10929), .Z(n9499) );
  MUX2_X2 U14090 ( .A(n9499), .B(n9492), .S(n10947), .Z(n9500) );
  MUX2_X2 U14091 ( .A(decode_regfile_intregs_14__22_), .B(
        decode_regfile_intregs_15__22_), .S(n10809), .Z(n9501) );
  MUX2_X2 U14092 ( .A(decode_regfile_intregs_12__22_), .B(
        decode_regfile_intregs_13__22_), .S(n10809), .Z(n9502) );
  MUX2_X2 U14093 ( .A(n9502), .B(n9501), .S(n10895), .Z(n9503) );
  MUX2_X2 U14094 ( .A(decode_regfile_intregs_10__22_), .B(
        decode_regfile_intregs_11__22_), .S(n10809), .Z(n9504) );
  MUX2_X2 U14095 ( .A(decode_regfile_intregs_8__22_), .B(
        decode_regfile_intregs_9__22_), .S(n10809), .Z(n9505) );
  MUX2_X2 U14096 ( .A(n9505), .B(n9504), .S(n10895), .Z(n9506) );
  MUX2_X2 U14097 ( .A(n9506), .B(n9503), .S(n10929), .Z(n9507) );
  MUX2_X2 U14098 ( .A(decode_regfile_intregs_6__22_), .B(
        decode_regfile_intregs_7__22_), .S(n10810), .Z(n9508) );
  MUX2_X2 U14099 ( .A(decode_regfile_intregs_4__22_), .B(
        decode_regfile_intregs_5__22_), .S(n10810), .Z(n9509) );
  MUX2_X2 U14100 ( .A(n9509), .B(n9508), .S(n10896), .Z(n9510) );
  MUX2_X2 U14101 ( .A(decode_regfile_intregs_2__22_), .B(
        decode_regfile_intregs_3__22_), .S(n10810), .Z(n9511) );
  MUX2_X2 U14102 ( .A(decode_regfile_intregs_0__22_), .B(
        decode_regfile_intregs_1__22_), .S(n10810), .Z(n9512) );
  MUX2_X2 U14103 ( .A(n9512), .B(n9511), .S(n10896), .Z(n9513) );
  MUX2_X2 U14104 ( .A(n9513), .B(n9510), .S(n10930), .Z(n9514) );
  MUX2_X2 U14105 ( .A(n9514), .B(n9507), .S(n10947), .Z(n9515) );
  MUX2_X2 U14106 ( .A(n9515), .B(n9500), .S(n10957), .Z(decode_regfile_N69) );
  MUX2_X2 U14107 ( .A(decode_regfile_intregs_30__23_), .B(
        decode_regfile_intregs_31__23_), .S(n10810), .Z(n9516) );
  MUX2_X2 U14108 ( .A(decode_regfile_intregs_28__23_), .B(
        decode_regfile_intregs_29__23_), .S(n10810), .Z(n9517) );
  MUX2_X2 U14109 ( .A(n9517), .B(n9516), .S(n10896), .Z(n9518) );
  MUX2_X2 U14110 ( .A(decode_regfile_intregs_26__23_), .B(
        decode_regfile_intregs_27__23_), .S(n10810), .Z(n9519) );
  MUX2_X2 U14111 ( .A(decode_regfile_intregs_24__23_), .B(
        decode_regfile_intregs_25__23_), .S(n10810), .Z(n9520) );
  MUX2_X2 U14112 ( .A(n9520), .B(n9519), .S(n10896), .Z(n9521) );
  MUX2_X2 U14113 ( .A(n9521), .B(n9518), .S(n10930), .Z(n9522) );
  MUX2_X2 U14114 ( .A(decode_regfile_intregs_22__23_), .B(
        decode_regfile_intregs_23__23_), .S(n10810), .Z(n9523) );
  MUX2_X2 U14115 ( .A(decode_regfile_intregs_20__23_), .B(
        decode_regfile_intregs_21__23_), .S(n10810), .Z(n9524) );
  MUX2_X2 U14116 ( .A(n9524), .B(n9523), .S(n10896), .Z(n9525) );
  MUX2_X2 U14117 ( .A(decode_regfile_intregs_18__23_), .B(
        decode_regfile_intregs_19__23_), .S(n10810), .Z(n9526) );
  MUX2_X2 U14118 ( .A(decode_regfile_intregs_16__23_), .B(
        decode_regfile_intregs_17__23_), .S(n10811), .Z(n9527) );
  MUX2_X2 U14119 ( .A(n9527), .B(n9526), .S(n10896), .Z(n9528) );
  MUX2_X2 U14120 ( .A(n9528), .B(n9525), .S(n10930), .Z(n9529) );
  MUX2_X2 U14121 ( .A(n9529), .B(n9522), .S(n10947), .Z(n9530) );
  MUX2_X2 U14122 ( .A(decode_regfile_intregs_14__23_), .B(
        decode_regfile_intregs_15__23_), .S(n10811), .Z(n9531) );
  MUX2_X2 U14123 ( .A(decode_regfile_intregs_12__23_), .B(
        decode_regfile_intregs_13__23_), .S(n10811), .Z(n9532) );
  MUX2_X2 U14124 ( .A(n9532), .B(n9531), .S(n10896), .Z(n9533) );
  MUX2_X2 U14125 ( .A(decode_regfile_intregs_10__23_), .B(
        decode_regfile_intregs_11__23_), .S(n10811), .Z(n9534) );
  MUX2_X2 U14126 ( .A(decode_regfile_intregs_8__23_), .B(
        decode_regfile_intregs_9__23_), .S(n10811), .Z(n9535) );
  MUX2_X2 U14127 ( .A(n9535), .B(n9534), .S(n10896), .Z(n9536) );
  MUX2_X2 U14128 ( .A(n9536), .B(n9533), .S(n10930), .Z(n9537) );
  MUX2_X2 U14129 ( .A(decode_regfile_intregs_6__23_), .B(
        decode_regfile_intregs_7__23_), .S(n10811), .Z(n9538) );
  MUX2_X2 U14130 ( .A(decode_regfile_intregs_4__23_), .B(
        decode_regfile_intregs_5__23_), .S(n10811), .Z(n9539) );
  MUX2_X2 U14131 ( .A(n9539), .B(n9538), .S(n10896), .Z(n9540) );
  MUX2_X2 U14132 ( .A(decode_regfile_intregs_2__23_), .B(
        decode_regfile_intregs_3__23_), .S(n10811), .Z(n9541) );
  MUX2_X2 U14133 ( .A(decode_regfile_intregs_0__23_), .B(
        decode_regfile_intregs_1__23_), .S(n10811), .Z(n9542) );
  MUX2_X2 U14134 ( .A(n9542), .B(n9541), .S(n10896), .Z(n9543) );
  MUX2_X2 U14135 ( .A(n9543), .B(n9540), .S(n10930), .Z(n9544) );
  MUX2_X2 U14136 ( .A(n9544), .B(n9537), .S(n10947), .Z(n9545) );
  MUX2_X2 U14137 ( .A(n9545), .B(n9530), .S(n10957), .Z(decode_regfile_N68) );
  MUX2_X2 U14138 ( .A(decode_regfile_intregs_30__24_), .B(
        decode_regfile_intregs_31__24_), .S(n10811), .Z(n9546) );
  MUX2_X2 U14139 ( .A(decode_regfile_intregs_28__24_), .B(
        decode_regfile_intregs_29__24_), .S(n10811), .Z(n9547) );
  MUX2_X2 U14140 ( .A(n9547), .B(n9546), .S(n10896), .Z(n9548) );
  MUX2_X2 U14141 ( .A(decode_regfile_intregs_26__24_), .B(
        decode_regfile_intregs_27__24_), .S(n10812), .Z(n9549) );
  MUX2_X2 U14142 ( .A(decode_regfile_intregs_24__24_), .B(
        decode_regfile_intregs_25__24_), .S(n10812), .Z(n9550) );
  MUX2_X2 U14143 ( .A(n9550), .B(n9549), .S(n10897), .Z(n9551) );
  MUX2_X2 U14144 ( .A(n9551), .B(n9548), .S(n10930), .Z(n9552) );
  MUX2_X2 U14145 ( .A(decode_regfile_intregs_22__24_), .B(
        decode_regfile_intregs_23__24_), .S(n10812), .Z(n9553) );
  MUX2_X2 U14146 ( .A(decode_regfile_intregs_20__24_), .B(
        decode_regfile_intregs_21__24_), .S(n10812), .Z(n9554) );
  MUX2_X2 U14147 ( .A(n9554), .B(n9553), .S(n10897), .Z(n9555) );
  MUX2_X2 U14148 ( .A(decode_regfile_intregs_18__24_), .B(
        decode_regfile_intregs_19__24_), .S(n10812), .Z(n9556) );
  MUX2_X2 U14149 ( .A(decode_regfile_intregs_16__24_), .B(
        decode_regfile_intregs_17__24_), .S(n10812), .Z(n9557) );
  MUX2_X2 U14150 ( .A(n9557), .B(n9556), .S(n10897), .Z(n9558) );
  MUX2_X2 U14151 ( .A(n9558), .B(n9555), .S(n10930), .Z(n9559) );
  MUX2_X2 U14152 ( .A(n9559), .B(n9552), .S(n10947), .Z(n9560) );
  MUX2_X2 U14153 ( .A(decode_regfile_intregs_14__24_), .B(
        decode_regfile_intregs_15__24_), .S(n10812), .Z(n9561) );
  MUX2_X2 U14154 ( .A(decode_regfile_intregs_12__24_), .B(
        decode_regfile_intregs_13__24_), .S(n10812), .Z(n9562) );
  MUX2_X2 U14155 ( .A(n9562), .B(n9561), .S(n10897), .Z(n9563) );
  MUX2_X2 U14156 ( .A(decode_regfile_intregs_10__24_), .B(
        decode_regfile_intregs_11__24_), .S(n10812), .Z(n9564) );
  MUX2_X2 U14157 ( .A(decode_regfile_intregs_8__24_), .B(
        decode_regfile_intregs_9__24_), .S(n10812), .Z(n9565) );
  MUX2_X2 U14158 ( .A(n9565), .B(n9564), .S(n10897), .Z(n9566) );
  MUX2_X2 U14159 ( .A(n9566), .B(n9563), .S(n10930), .Z(n9567) );
  MUX2_X2 U14160 ( .A(decode_regfile_intregs_6__24_), .B(
        decode_regfile_intregs_7__24_), .S(n10812), .Z(n9568) );
  MUX2_X2 U14161 ( .A(decode_regfile_intregs_4__24_), .B(
        decode_regfile_intregs_5__24_), .S(n10813), .Z(n9569) );
  MUX2_X2 U14162 ( .A(n9569), .B(n9568), .S(n10897), .Z(n9570) );
  MUX2_X2 U14163 ( .A(decode_regfile_intregs_2__24_), .B(
        decode_regfile_intregs_3__24_), .S(n10813), .Z(n9571) );
  MUX2_X2 U14164 ( .A(decode_regfile_intregs_0__24_), .B(
        decode_regfile_intregs_1__24_), .S(n10813), .Z(n9572) );
  MUX2_X2 U14165 ( .A(n9572), .B(n9571), .S(n10897), .Z(n9573) );
  MUX2_X2 U14166 ( .A(n9573), .B(n9570), .S(n10930), .Z(n9574) );
  MUX2_X2 U14167 ( .A(n9574), .B(n9567), .S(n10947), .Z(n9575) );
  MUX2_X2 U14168 ( .A(n9575), .B(n9560), .S(n10957), .Z(decode_regfile_N67) );
  MUX2_X2 U14169 ( .A(decode_regfile_intregs_30__25_), .B(
        decode_regfile_intregs_31__25_), .S(n10813), .Z(n9576) );
  MUX2_X2 U14170 ( .A(decode_regfile_intregs_28__25_), .B(
        decode_regfile_intregs_29__25_), .S(n10813), .Z(n9577) );
  MUX2_X2 U14171 ( .A(n9577), .B(n9576), .S(n10897), .Z(n9578) );
  MUX2_X2 U14172 ( .A(decode_regfile_intregs_26__25_), .B(
        decode_regfile_intregs_27__25_), .S(n10813), .Z(n9579) );
  MUX2_X2 U14173 ( .A(decode_regfile_intregs_24__25_), .B(
        decode_regfile_intregs_25__25_), .S(n10813), .Z(n9580) );
  MUX2_X2 U14174 ( .A(n9580), .B(n9579), .S(n10897), .Z(n9581) );
  MUX2_X2 U14175 ( .A(n9581), .B(n9578), .S(n10930), .Z(n9582) );
  MUX2_X2 U14176 ( .A(decode_regfile_intregs_22__25_), .B(
        decode_regfile_intregs_23__25_), .S(n10813), .Z(n9583) );
  MUX2_X2 U14177 ( .A(decode_regfile_intregs_20__25_), .B(
        decode_regfile_intregs_21__25_), .S(n10813), .Z(n9584) );
  MUX2_X2 U14178 ( .A(n9584), .B(n9583), .S(n10897), .Z(n9585) );
  MUX2_X2 U14179 ( .A(decode_regfile_intregs_18__25_), .B(
        decode_regfile_intregs_19__25_), .S(n10813), .Z(n9586) );
  MUX2_X2 U14180 ( .A(decode_regfile_intregs_16__25_), .B(
        decode_regfile_intregs_17__25_), .S(n10813), .Z(n9587) );
  MUX2_X2 U14181 ( .A(n9587), .B(n9586), .S(n10897), .Z(n9588) );
  MUX2_X2 U14182 ( .A(n9588), .B(n9585), .S(n10930), .Z(n9589) );
  MUX2_X2 U14183 ( .A(n9589), .B(n9582), .S(n10947), .Z(n9590) );
  MUX2_X2 U14184 ( .A(decode_regfile_intregs_14__25_), .B(
        decode_regfile_intregs_15__25_), .S(n10814), .Z(n9591) );
  MUX2_X2 U14185 ( .A(decode_regfile_intregs_12__25_), .B(
        decode_regfile_intregs_13__25_), .S(n10814), .Z(n9592) );
  MUX2_X2 U14186 ( .A(n9592), .B(n9591), .S(n10898), .Z(n9593) );
  MUX2_X2 U14187 ( .A(decode_regfile_intregs_10__25_), .B(
        decode_regfile_intregs_11__25_), .S(n10814), .Z(n9594) );
  MUX2_X2 U14188 ( .A(decode_regfile_intregs_8__25_), .B(
        decode_regfile_intregs_9__25_), .S(n10814), .Z(n9595) );
  MUX2_X2 U14189 ( .A(n9595), .B(n9594), .S(n10898), .Z(n9596) );
  MUX2_X2 U14190 ( .A(n9596), .B(n9593), .S(n10931), .Z(n9597) );
  MUX2_X2 U14191 ( .A(decode_regfile_intregs_6__25_), .B(
        decode_regfile_intregs_7__25_), .S(n10814), .Z(n9598) );
  MUX2_X2 U14192 ( .A(decode_regfile_intregs_4__25_), .B(
        decode_regfile_intregs_5__25_), .S(n10814), .Z(n9599) );
  MUX2_X2 U14193 ( .A(n9599), .B(n9598), .S(n10898), .Z(n9600) );
  MUX2_X2 U14194 ( .A(decode_regfile_intregs_2__25_), .B(
        decode_regfile_intregs_3__25_), .S(n10814), .Z(n9601) );
  MUX2_X2 U14195 ( .A(decode_regfile_intregs_0__25_), .B(
        decode_regfile_intregs_1__25_), .S(n10814), .Z(n9602) );
  MUX2_X2 U14196 ( .A(n9602), .B(n9601), .S(n10898), .Z(n9603) );
  MUX2_X2 U14197 ( .A(n9603), .B(n9600), .S(n10931), .Z(n9604) );
  MUX2_X2 U14198 ( .A(n9604), .B(n9597), .S(n10948), .Z(n9605) );
  MUX2_X2 U14199 ( .A(n9605), .B(n9590), .S(n10957), .Z(decode_regfile_N66) );
  MUX2_X2 U14200 ( .A(decode_regfile_intregs_30__26_), .B(
        decode_regfile_intregs_31__26_), .S(n10814), .Z(n9606) );
  MUX2_X2 U14201 ( .A(decode_regfile_intregs_28__26_), .B(
        decode_regfile_intregs_29__26_), .S(n10814), .Z(n9607) );
  MUX2_X2 U14202 ( .A(n9607), .B(n9606), .S(n10898), .Z(n9608) );
  MUX2_X2 U14203 ( .A(decode_regfile_intregs_26__26_), .B(
        decode_regfile_intregs_27__26_), .S(n10814), .Z(n9609) );
  MUX2_X2 U14204 ( .A(decode_regfile_intregs_24__26_), .B(
        decode_regfile_intregs_25__26_), .S(n10815), .Z(n9610) );
  MUX2_X2 U14205 ( .A(n9610), .B(n9609), .S(n10898), .Z(n9611) );
  MUX2_X2 U14206 ( .A(n9611), .B(n9608), .S(n10931), .Z(n9612) );
  MUX2_X2 U14207 ( .A(decode_regfile_intregs_22__26_), .B(
        decode_regfile_intregs_23__26_), .S(n10815), .Z(n9613) );
  MUX2_X2 U14208 ( .A(decode_regfile_intregs_20__26_), .B(
        decode_regfile_intregs_21__26_), .S(n10815), .Z(n9614) );
  MUX2_X2 U14209 ( .A(n9614), .B(n9613), .S(n10898), .Z(n9615) );
  MUX2_X2 U14210 ( .A(decode_regfile_intregs_18__26_), .B(
        decode_regfile_intregs_19__26_), .S(n10815), .Z(n9616) );
  MUX2_X2 U14211 ( .A(decode_regfile_intregs_16__26_), .B(
        decode_regfile_intregs_17__26_), .S(n10815), .Z(n9617) );
  MUX2_X2 U14212 ( .A(n9617), .B(n9616), .S(n10898), .Z(n9618) );
  MUX2_X2 U14213 ( .A(n9618), .B(n9615), .S(n10931), .Z(n9619) );
  MUX2_X2 U14214 ( .A(n9619), .B(n9612), .S(n10948), .Z(n9620) );
  MUX2_X2 U14215 ( .A(decode_regfile_intregs_14__26_), .B(
        decode_regfile_intregs_15__26_), .S(n10815), .Z(n9621) );
  MUX2_X2 U14216 ( .A(decode_regfile_intregs_12__26_), .B(
        decode_regfile_intregs_13__26_), .S(n10815), .Z(n9622) );
  MUX2_X2 U14217 ( .A(n9622), .B(n9621), .S(n10898), .Z(n9623) );
  MUX2_X2 U14218 ( .A(decode_regfile_intregs_10__26_), .B(
        decode_regfile_intregs_11__26_), .S(n10815), .Z(n9624) );
  MUX2_X2 U14219 ( .A(decode_regfile_intregs_8__26_), .B(
        decode_regfile_intregs_9__26_), .S(n10815), .Z(n9625) );
  MUX2_X2 U14220 ( .A(n9625), .B(n9624), .S(n10898), .Z(n9626) );
  MUX2_X2 U14221 ( .A(n9626), .B(n9623), .S(n10931), .Z(n9627) );
  MUX2_X2 U14222 ( .A(decode_regfile_intregs_6__26_), .B(
        decode_regfile_intregs_7__26_), .S(n10815), .Z(n9628) );
  MUX2_X2 U14223 ( .A(decode_regfile_intregs_4__26_), .B(
        decode_regfile_intregs_5__26_), .S(n10815), .Z(n9629) );
  MUX2_X2 U14224 ( .A(n9629), .B(n9628), .S(n10898), .Z(n9630) );
  MUX2_X2 U14225 ( .A(decode_regfile_intregs_2__26_), .B(
        decode_regfile_intregs_3__26_), .S(n10816), .Z(n9631) );
  MUX2_X2 U14226 ( .A(decode_regfile_intregs_0__26_), .B(
        decode_regfile_intregs_1__26_), .S(n10816), .Z(n9632) );
  MUX2_X2 U14227 ( .A(n9632), .B(n9631), .S(n10899), .Z(n9633) );
  MUX2_X2 U14228 ( .A(n9633), .B(n9630), .S(n10931), .Z(n9634) );
  MUX2_X2 U14229 ( .A(n9634), .B(n9627), .S(n10948), .Z(n9635) );
  MUX2_X2 U14230 ( .A(n9635), .B(n9620), .S(n10957), .Z(decode_regfile_N65) );
  MUX2_X2 U14231 ( .A(decode_regfile_intregs_30__27_), .B(
        decode_regfile_intregs_31__27_), .S(n10816), .Z(n9636) );
  MUX2_X2 U14232 ( .A(decode_regfile_intregs_28__27_), .B(
        decode_regfile_intregs_29__27_), .S(n10816), .Z(n9637) );
  MUX2_X2 U14233 ( .A(n9637), .B(n9636), .S(n10899), .Z(n9638) );
  MUX2_X2 U14234 ( .A(decode_regfile_intregs_26__27_), .B(
        decode_regfile_intregs_27__27_), .S(n10816), .Z(n9639) );
  MUX2_X2 U14235 ( .A(decode_regfile_intregs_24__27_), .B(
        decode_regfile_intregs_25__27_), .S(n10816), .Z(n9640) );
  MUX2_X2 U14236 ( .A(n9640), .B(n9639), .S(n10899), .Z(n9641) );
  MUX2_X2 U14237 ( .A(n9641), .B(n9638), .S(n10931), .Z(n9642) );
  MUX2_X2 U14238 ( .A(decode_regfile_intregs_22__27_), .B(
        decode_regfile_intregs_23__27_), .S(n10816), .Z(n9643) );
  MUX2_X2 U14239 ( .A(decode_regfile_intregs_20__27_), .B(
        decode_regfile_intregs_21__27_), .S(n10816), .Z(n9644) );
  MUX2_X2 U14240 ( .A(n9644), .B(n9643), .S(n10899), .Z(n9645) );
  MUX2_X2 U14241 ( .A(decode_regfile_intregs_18__27_), .B(
        decode_regfile_intregs_19__27_), .S(n10816), .Z(n9646) );
  MUX2_X2 U14242 ( .A(decode_regfile_intregs_16__27_), .B(
        decode_regfile_intregs_17__27_), .S(n10816), .Z(n9647) );
  MUX2_X2 U14243 ( .A(n9647), .B(n9646), .S(n10899), .Z(n9648) );
  MUX2_X2 U14244 ( .A(n9648), .B(n9645), .S(n10931), .Z(n9649) );
  MUX2_X2 U14245 ( .A(n9649), .B(n9642), .S(n10948), .Z(n9650) );
  MUX2_X2 U14246 ( .A(decode_regfile_intregs_14__27_), .B(
        decode_regfile_intregs_15__27_), .S(n10816), .Z(n9651) );
  MUX2_X2 U14247 ( .A(decode_regfile_intregs_12__27_), .B(
        decode_regfile_intregs_13__27_), .S(n10817), .Z(n9652) );
  MUX2_X2 U14248 ( .A(n9652), .B(n9651), .S(n10899), .Z(n9653) );
  MUX2_X2 U14249 ( .A(decode_regfile_intregs_10__27_), .B(
        decode_regfile_intregs_11__27_), .S(n10817), .Z(n9654) );
  MUX2_X2 U14250 ( .A(decode_regfile_intregs_8__27_), .B(
        decode_regfile_intregs_9__27_), .S(n10817), .Z(n9655) );
  MUX2_X2 U14251 ( .A(n9655), .B(n9654), .S(n10899), .Z(n9656) );
  MUX2_X2 U14252 ( .A(n9656), .B(n9653), .S(n10931), .Z(n9657) );
  MUX2_X2 U14253 ( .A(decode_regfile_intregs_6__27_), .B(
        decode_regfile_intregs_7__27_), .S(n10817), .Z(n9658) );
  MUX2_X2 U14254 ( .A(decode_regfile_intregs_4__27_), .B(
        decode_regfile_intregs_5__27_), .S(n10817), .Z(n9659) );
  MUX2_X2 U14255 ( .A(n9659), .B(n9658), .S(n10899), .Z(n9660) );
  MUX2_X2 U14256 ( .A(decode_regfile_intregs_2__27_), .B(
        decode_regfile_intregs_3__27_), .S(n10817), .Z(n9661) );
  MUX2_X2 U14257 ( .A(decode_regfile_intregs_0__27_), .B(
        decode_regfile_intregs_1__27_), .S(n10817), .Z(n9662) );
  MUX2_X2 U14258 ( .A(n9662), .B(n9661), .S(n10899), .Z(n9663) );
  MUX2_X2 U14259 ( .A(n9663), .B(n9660), .S(n10931), .Z(n9664) );
  MUX2_X2 U14260 ( .A(n9664), .B(n9657), .S(n10948), .Z(n9665) );
  MUX2_X2 U14261 ( .A(n9665), .B(n9650), .S(n10957), .Z(decode_regfile_N64) );
  MUX2_X2 U14262 ( .A(decode_regfile_intregs_30__28_), .B(
        decode_regfile_intregs_31__28_), .S(n10817), .Z(n9666) );
  MUX2_X2 U14263 ( .A(decode_regfile_intregs_28__28_), .B(
        decode_regfile_intregs_29__28_), .S(n10817), .Z(n9667) );
  MUX2_X2 U14264 ( .A(n9667), .B(n9666), .S(n10899), .Z(n9668) );
  MUX2_X2 U14265 ( .A(decode_regfile_intregs_26__28_), .B(
        decode_regfile_intregs_27__28_), .S(n10817), .Z(n9669) );
  MUX2_X2 U14266 ( .A(decode_regfile_intregs_24__28_), .B(
        decode_regfile_intregs_25__28_), .S(n10817), .Z(n9670) );
  MUX2_X2 U14267 ( .A(n9670), .B(n9669), .S(n10899), .Z(n9671) );
  MUX2_X2 U14268 ( .A(n9671), .B(n9668), .S(n10931), .Z(n9672) );
  MUX2_X2 U14269 ( .A(decode_regfile_intregs_22__28_), .B(
        decode_regfile_intregs_23__28_), .S(n10818), .Z(n9673) );
  MUX2_X2 U14270 ( .A(decode_regfile_intregs_20__28_), .B(
        decode_regfile_intregs_21__28_), .S(n10818), .Z(n9674) );
  MUX2_X2 U14271 ( .A(n9674), .B(n9673), .S(n10900), .Z(n9675) );
  MUX2_X2 U14272 ( .A(decode_regfile_intregs_18__28_), .B(
        decode_regfile_intregs_19__28_), .S(n10818), .Z(n9676) );
  MUX2_X2 U14273 ( .A(decode_regfile_intregs_16__28_), .B(
        decode_regfile_intregs_17__28_), .S(n10818), .Z(n9677) );
  MUX2_X2 U14274 ( .A(n9677), .B(n9676), .S(n10900), .Z(n9678) );
  MUX2_X2 U14275 ( .A(n9678), .B(n9675), .S(n10932), .Z(n9679) );
  MUX2_X2 U14276 ( .A(n9679), .B(n9672), .S(n10948), .Z(n9680) );
  MUX2_X2 U14277 ( .A(decode_regfile_intregs_14__28_), .B(
        decode_regfile_intregs_15__28_), .S(n10818), .Z(n9681) );
  MUX2_X2 U14278 ( .A(decode_regfile_intregs_12__28_), .B(
        decode_regfile_intregs_13__28_), .S(n10818), .Z(n9682) );
  MUX2_X2 U14279 ( .A(n9682), .B(n9681), .S(n10900), .Z(n9683) );
  MUX2_X2 U14280 ( .A(decode_regfile_intregs_10__28_), .B(
        decode_regfile_intregs_11__28_), .S(n10818), .Z(n9684) );
  MUX2_X2 U14281 ( .A(decode_regfile_intregs_8__28_), .B(
        decode_regfile_intregs_9__28_), .S(n10818), .Z(n9685) );
  MUX2_X2 U14282 ( .A(n9685), .B(n9684), .S(n10900), .Z(n9686) );
  MUX2_X2 U14283 ( .A(n9686), .B(n9683), .S(n10932), .Z(n9687) );
  MUX2_X2 U14284 ( .A(decode_regfile_intregs_6__28_), .B(
        decode_regfile_intregs_7__28_), .S(n10818), .Z(n9688) );
  MUX2_X2 U14285 ( .A(decode_regfile_intregs_4__28_), .B(
        decode_regfile_intregs_5__28_), .S(n10818), .Z(n9689) );
  MUX2_X2 U14286 ( .A(n9689), .B(n9688), .S(n10900), .Z(n9690) );
  MUX2_X2 U14287 ( .A(decode_regfile_intregs_2__28_), .B(
        decode_regfile_intregs_3__28_), .S(n10818), .Z(n9691) );
  MUX2_X2 U14288 ( .A(decode_regfile_intregs_0__28_), .B(
        decode_regfile_intregs_1__28_), .S(n10819), .Z(n9692) );
  MUX2_X2 U14289 ( .A(n9692), .B(n9691), .S(n10900), .Z(n9693) );
  MUX2_X2 U14290 ( .A(n9693), .B(n9690), .S(n10932), .Z(n9694) );
  MUX2_X2 U14291 ( .A(n9694), .B(n9687), .S(n10948), .Z(n9695) );
  MUX2_X2 U14292 ( .A(n9695), .B(n9680), .S(n10957), .Z(decode_regfile_N63) );
  MUX2_X2 U14293 ( .A(decode_regfile_intregs_30__29_), .B(
        decode_regfile_intregs_31__29_), .S(n10819), .Z(n9696) );
  MUX2_X2 U14294 ( .A(decode_regfile_intregs_28__29_), .B(
        decode_regfile_intregs_29__29_), .S(n10819), .Z(n9697) );
  MUX2_X2 U14295 ( .A(n9697), .B(n9696), .S(n10900), .Z(n9698) );
  MUX2_X2 U14296 ( .A(decode_regfile_intregs_26__29_), .B(
        decode_regfile_intregs_27__29_), .S(n10819), .Z(n9699) );
  MUX2_X2 U14297 ( .A(decode_regfile_intregs_24__29_), .B(
        decode_regfile_intregs_25__29_), .S(n10819), .Z(n9700) );
  MUX2_X2 U14298 ( .A(n9700), .B(n9699), .S(n10900), .Z(n9701) );
  MUX2_X2 U14299 ( .A(n9701), .B(n9698), .S(n10932), .Z(n9702) );
  MUX2_X2 U14300 ( .A(decode_regfile_intregs_22__29_), .B(
        decode_regfile_intregs_23__29_), .S(n10819), .Z(n9703) );
  MUX2_X2 U14301 ( .A(decode_regfile_intregs_20__29_), .B(
        decode_regfile_intregs_21__29_), .S(n10819), .Z(n9704) );
  MUX2_X2 U14302 ( .A(n9704), .B(n9703), .S(n10900), .Z(n9705) );
  MUX2_X2 U14303 ( .A(decode_regfile_intregs_18__29_), .B(
        decode_regfile_intregs_19__29_), .S(n10819), .Z(n9706) );
  MUX2_X2 U14304 ( .A(decode_regfile_intregs_16__29_), .B(
        decode_regfile_intregs_17__29_), .S(n10819), .Z(n9707) );
  MUX2_X2 U14305 ( .A(n9707), .B(n9706), .S(n10900), .Z(n9708) );
  MUX2_X2 U14306 ( .A(n9708), .B(n9705), .S(n10932), .Z(n9709) );
  MUX2_X2 U14307 ( .A(n9709), .B(n9702), .S(n10948), .Z(n9710) );
  MUX2_X2 U14308 ( .A(decode_regfile_intregs_14__29_), .B(
        decode_regfile_intregs_15__29_), .S(n10819), .Z(n9711) );
  MUX2_X2 U14309 ( .A(decode_regfile_intregs_12__29_), .B(
        decode_regfile_intregs_13__29_), .S(n10819), .Z(n9712) );
  MUX2_X2 U14310 ( .A(n9712), .B(n9711), .S(n10900), .Z(n9713) );
  MUX2_X2 U14311 ( .A(decode_regfile_intregs_10__29_), .B(
        decode_regfile_intregs_11__29_), .S(n10820), .Z(n9714) );
  MUX2_X2 U14312 ( .A(decode_regfile_intregs_8__29_), .B(
        decode_regfile_intregs_9__29_), .S(n10820), .Z(n9715) );
  MUX2_X2 U14313 ( .A(n9715), .B(n9714), .S(n10901), .Z(n9716) );
  MUX2_X2 U14314 ( .A(n9716), .B(n9713), .S(n10932), .Z(n9717) );
  MUX2_X2 U14315 ( .A(decode_regfile_intregs_6__29_), .B(
        decode_regfile_intregs_7__29_), .S(n10820), .Z(n9718) );
  MUX2_X2 U14316 ( .A(decode_regfile_intregs_4__29_), .B(
        decode_regfile_intregs_5__29_), .S(n10820), .Z(n9719) );
  MUX2_X2 U14317 ( .A(n9719), .B(n9718), .S(n10901), .Z(n9720) );
  MUX2_X2 U14318 ( .A(decode_regfile_intregs_2__29_), .B(
        decode_regfile_intregs_3__29_), .S(n10820), .Z(n9721) );
  MUX2_X2 U14319 ( .A(decode_regfile_intregs_0__29_), .B(
        decode_regfile_intregs_1__29_), .S(n10820), .Z(n9722) );
  MUX2_X2 U14320 ( .A(n9722), .B(n9721), .S(n10901), .Z(n9723) );
  MUX2_X2 U14321 ( .A(n9723), .B(n9720), .S(n10932), .Z(n9724) );
  MUX2_X2 U14322 ( .A(n9724), .B(n9717), .S(n10948), .Z(n9725) );
  MUX2_X2 U14323 ( .A(n9725), .B(n9710), .S(n10957), .Z(decode_regfile_N62) );
  MUX2_X2 U14324 ( .A(decode_regfile_intregs_30__30_), .B(
        decode_regfile_intregs_31__30_), .S(n10820), .Z(n9726) );
  MUX2_X2 U14325 ( .A(decode_regfile_intregs_28__30_), .B(
        decode_regfile_intregs_29__30_), .S(n10820), .Z(n9727) );
  MUX2_X2 U14326 ( .A(n9727), .B(n9726), .S(n10901), .Z(n9728) );
  MUX2_X2 U14327 ( .A(decode_regfile_intregs_26__30_), .B(
        decode_regfile_intregs_27__30_), .S(n10820), .Z(n9729) );
  MUX2_X2 U14328 ( .A(decode_regfile_intregs_24__30_), .B(
        decode_regfile_intregs_25__30_), .S(n10820), .Z(n9730) );
  MUX2_X2 U14329 ( .A(n9730), .B(n9729), .S(n10901), .Z(n9731) );
  MUX2_X2 U14330 ( .A(n9731), .B(n9728), .S(n10932), .Z(n9732) );
  MUX2_X2 U14331 ( .A(decode_regfile_intregs_22__30_), .B(
        decode_regfile_intregs_23__30_), .S(n10820), .Z(n9733) );
  MUX2_X2 U14332 ( .A(decode_regfile_intregs_20__30_), .B(
        decode_regfile_intregs_21__30_), .S(n10821), .Z(n9734) );
  MUX2_X2 U14333 ( .A(n9734), .B(n9733), .S(n10901), .Z(n9735) );
  MUX2_X2 U14334 ( .A(decode_regfile_intregs_18__30_), .B(
        decode_regfile_intregs_19__30_), .S(n10821), .Z(n9736) );
  MUX2_X2 U14335 ( .A(decode_regfile_intregs_16__30_), .B(
        decode_regfile_intregs_17__30_), .S(n10821), .Z(n9737) );
  MUX2_X2 U14336 ( .A(n9737), .B(n9736), .S(n10901), .Z(n9738) );
  MUX2_X2 U14337 ( .A(n9738), .B(n9735), .S(n10932), .Z(n9739) );
  MUX2_X2 U14338 ( .A(n9739), .B(n9732), .S(n10948), .Z(n9740) );
  MUX2_X2 U14339 ( .A(decode_regfile_intregs_14__30_), .B(
        decode_regfile_intregs_15__30_), .S(n10821), .Z(n9741) );
  MUX2_X2 U14340 ( .A(decode_regfile_intregs_12__30_), .B(
        decode_regfile_intregs_13__30_), .S(n10821), .Z(n9742) );
  MUX2_X2 U14341 ( .A(n9742), .B(n9741), .S(n10901), .Z(n9743) );
  MUX2_X2 U14342 ( .A(decode_regfile_intregs_10__30_), .B(
        decode_regfile_intregs_11__30_), .S(n10821), .Z(n9744) );
  MUX2_X2 U14343 ( .A(decode_regfile_intregs_8__30_), .B(
        decode_regfile_intregs_9__30_), .S(n10821), .Z(n9745) );
  MUX2_X2 U14344 ( .A(n9745), .B(n9744), .S(n10901), .Z(n9746) );
  MUX2_X2 U14345 ( .A(n9746), .B(n9743), .S(n10932), .Z(n9747) );
  MUX2_X2 U14346 ( .A(decode_regfile_intregs_6__30_), .B(
        decode_regfile_intregs_7__30_), .S(n10821), .Z(n9748) );
  MUX2_X2 U14347 ( .A(decode_regfile_intregs_4__30_), .B(
        decode_regfile_intregs_5__30_), .S(n10821), .Z(n9749) );
  MUX2_X2 U14348 ( .A(n9749), .B(n9748), .S(n10901), .Z(n9750) );
  MUX2_X2 U14349 ( .A(decode_regfile_intregs_2__30_), .B(
        decode_regfile_intregs_3__30_), .S(n10821), .Z(n9751) );
  MUX2_X2 U14350 ( .A(decode_regfile_intregs_0__30_), .B(
        decode_regfile_intregs_1__30_), .S(n10821), .Z(n9752) );
  MUX2_X2 U14351 ( .A(n9752), .B(n9751), .S(n10901), .Z(n9753) );
  MUX2_X2 U14352 ( .A(n9753), .B(n9750), .S(n10932), .Z(n9754) );
  MUX2_X2 U14353 ( .A(n9754), .B(n9747), .S(n10948), .Z(n9755) );
  MUX2_X2 U14354 ( .A(n9755), .B(n9740), .S(n10957), .Z(decode_regfile_N61) );
  MUX2_X2 U14355 ( .A(decode_regfile_intregs_30__31_), .B(
        decode_regfile_intregs_31__31_), .S(n10822), .Z(n9756) );
  MUX2_X2 U14356 ( .A(decode_regfile_intregs_28__31_), .B(
        decode_regfile_intregs_29__31_), .S(n10822), .Z(n9757) );
  MUX2_X2 U14357 ( .A(n9757), .B(n9756), .S(n10902), .Z(n9758) );
  MUX2_X2 U14358 ( .A(decode_regfile_intregs_26__31_), .B(
        decode_regfile_intregs_27__31_), .S(n10822), .Z(n9759) );
  MUX2_X2 U14359 ( .A(decode_regfile_intregs_24__31_), .B(
        decode_regfile_intregs_25__31_), .S(n10822), .Z(n9760) );
  MUX2_X2 U14360 ( .A(n9760), .B(n9759), .S(n10902), .Z(n9761) );
  MUX2_X2 U14361 ( .A(n9761), .B(n9758), .S(n10933), .Z(n9762) );
  MUX2_X2 U14362 ( .A(decode_regfile_intregs_22__31_), .B(
        decode_regfile_intregs_23__31_), .S(n10822), .Z(n9763) );
  MUX2_X2 U14363 ( .A(decode_regfile_intregs_20__31_), .B(
        decode_regfile_intregs_21__31_), .S(n10822), .Z(n9764) );
  MUX2_X2 U14364 ( .A(n9764), .B(n9763), .S(n10902), .Z(n9765) );
  MUX2_X2 U14365 ( .A(decode_regfile_intregs_18__31_), .B(
        decode_regfile_intregs_19__31_), .S(n10822), .Z(n9766) );
  MUX2_X2 U14366 ( .A(decode_regfile_intregs_16__31_), .B(
        decode_regfile_intregs_17__31_), .S(n10822), .Z(n9767) );
  MUX2_X2 U14367 ( .A(n9767), .B(n9766), .S(n10902), .Z(n9768) );
  MUX2_X2 U14368 ( .A(n9768), .B(n9765), .S(n10933), .Z(n9769) );
  MUX2_X2 U14369 ( .A(n9769), .B(n9762), .S(n10949), .Z(n9770) );
  MUX2_X2 U14370 ( .A(decode_regfile_intregs_14__31_), .B(
        decode_regfile_intregs_15__31_), .S(n10822), .Z(n9771) );
  MUX2_X2 U14371 ( .A(decode_regfile_intregs_12__31_), .B(
        decode_regfile_intregs_13__31_), .S(n10822), .Z(n9772) );
  MUX2_X2 U14372 ( .A(n9772), .B(n9771), .S(n10902), .Z(n9773) );
  MUX2_X2 U14373 ( .A(decode_regfile_intregs_10__31_), .B(
        decode_regfile_intregs_11__31_), .S(n10822), .Z(n9774) );
  MUX2_X2 U14374 ( .A(decode_regfile_intregs_8__31_), .B(
        decode_regfile_intregs_9__31_), .S(n10823), .Z(n9775) );
  MUX2_X2 U14375 ( .A(n9775), .B(n9774), .S(n10902), .Z(n9776) );
  MUX2_X2 U14376 ( .A(n9776), .B(n9773), .S(n10933), .Z(n9777) );
  MUX2_X2 U14377 ( .A(decode_regfile_intregs_6__31_), .B(
        decode_regfile_intregs_7__31_), .S(n10823), .Z(n9778) );
  MUX2_X2 U14378 ( .A(decode_regfile_intregs_4__31_), .B(
        decode_regfile_intregs_5__31_), .S(n10823), .Z(n9779) );
  MUX2_X2 U14379 ( .A(n9779), .B(n9778), .S(n10902), .Z(n9780) );
  MUX2_X2 U14380 ( .A(decode_regfile_intregs_2__31_), .B(
        decode_regfile_intregs_3__31_), .S(n10823), .Z(n9781) );
  MUX2_X2 U14381 ( .A(decode_regfile_intregs_0__31_), .B(
        decode_regfile_intregs_1__31_), .S(n10823), .Z(n9782) );
  MUX2_X2 U14382 ( .A(n9782), .B(n9781), .S(n10902), .Z(n9783) );
  MUX2_X2 U14383 ( .A(n9783), .B(n9780), .S(n10933), .Z(n9784) );
  MUX2_X2 U14384 ( .A(n9784), .B(n9777), .S(n10949), .Z(n9785) );
  MUX2_X2 U14385 ( .A(n9785), .B(n9770), .S(n10958), .Z(decode_regfile_N60) );
  MUX2_X2 U14386 ( .A(decode_regfile_fpregs_30__0_), .B(
        decode_regfile_fpregs_31__0_), .S(n10823), .Z(n9786) );
  MUX2_X2 U14387 ( .A(decode_regfile_fpregs_28__0_), .B(
        decode_regfile_fpregs_29__0_), .S(n10823), .Z(n9787) );
  MUX2_X2 U14388 ( .A(n9787), .B(n9786), .S(n10902), .Z(n9788) );
  MUX2_X2 U14389 ( .A(decode_regfile_fpregs_26__0_), .B(
        decode_regfile_fpregs_27__0_), .S(n10823), .Z(n9789) );
  MUX2_X2 U14390 ( .A(decode_regfile_fpregs_24__0_), .B(
        decode_regfile_fpregs_25__0_), .S(n10823), .Z(n9790) );
  MUX2_X2 U14391 ( .A(n9790), .B(n9789), .S(n10902), .Z(n9791) );
  MUX2_X2 U14392 ( .A(n9791), .B(n9788), .S(n10933), .Z(n9792) );
  MUX2_X2 U14393 ( .A(decode_regfile_fpregs_22__0_), .B(
        decode_regfile_fpregs_23__0_), .S(n10823), .Z(n9793) );
  MUX2_X2 U14394 ( .A(decode_regfile_fpregs_20__0_), .B(
        decode_regfile_fpregs_21__0_), .S(n10823), .Z(n9794) );
  MUX2_X2 U14395 ( .A(n9794), .B(n9793), .S(n10902), .Z(n9795) );
  MUX2_X2 U14396 ( .A(decode_regfile_fpregs_18__0_), .B(
        decode_regfile_fpregs_19__0_), .S(n10824), .Z(n9796) );
  MUX2_X2 U14397 ( .A(decode_regfile_fpregs_16__0_), .B(
        decode_regfile_fpregs_17__0_), .S(n10824), .Z(n9797) );
  MUX2_X2 U14398 ( .A(n9797), .B(n9796), .S(n10903), .Z(n9798) );
  MUX2_X2 U14399 ( .A(n9798), .B(n9795), .S(n10933), .Z(n9799) );
  MUX2_X2 U14400 ( .A(n9799), .B(n9792), .S(n10949), .Z(n9800) );
  MUX2_X2 U14401 ( .A(decode_regfile_fpregs_14__0_), .B(
        decode_regfile_fpregs_15__0_), .S(n10824), .Z(n9801) );
  MUX2_X2 U14402 ( .A(decode_regfile_fpregs_12__0_), .B(
        decode_regfile_fpregs_13__0_), .S(n10824), .Z(n9802) );
  MUX2_X2 U14403 ( .A(n9802), .B(n9801), .S(n10903), .Z(n9803) );
  MUX2_X2 U14404 ( .A(decode_regfile_fpregs_10__0_), .B(
        decode_regfile_fpregs_11__0_), .S(n10824), .Z(n9804) );
  MUX2_X2 U14405 ( .A(decode_regfile_fpregs_8__0_), .B(
        decode_regfile_fpregs_9__0_), .S(n10824), .Z(n9805) );
  MUX2_X2 U14406 ( .A(n9805), .B(n9804), .S(n10903), .Z(n9806) );
  MUX2_X2 U14407 ( .A(n9806), .B(n9803), .S(n10933), .Z(n9807) );
  MUX2_X2 U14408 ( .A(decode_regfile_fpregs_6__0_), .B(
        decode_regfile_fpregs_7__0_), .S(n10824), .Z(n9808) );
  MUX2_X2 U14409 ( .A(decode_regfile_fpregs_4__0_), .B(
        decode_regfile_fpregs_5__0_), .S(n10824), .Z(n9809) );
  MUX2_X2 U14410 ( .A(n9809), .B(n9808), .S(n10903), .Z(n9810) );
  MUX2_X2 U14411 ( .A(decode_regfile_fpregs_2__0_), .B(
        decode_regfile_fpregs_3__0_), .S(n10824), .Z(n9811) );
  MUX2_X2 U14412 ( .A(decode_regfile_fpregs_0__0_), .B(
        decode_regfile_fpregs_1__0_), .S(n10824), .Z(n9812) );
  MUX2_X2 U14413 ( .A(n9812), .B(n9811), .S(n10903), .Z(n9813) );
  MUX2_X2 U14414 ( .A(n9813), .B(n9810), .S(n10933), .Z(n9814) );
  MUX2_X2 U14415 ( .A(n9814), .B(n9807), .S(n10949), .Z(n9815) );
  MUX2_X2 U14416 ( .A(n9815), .B(n9800), .S(n10958), .Z(decode_regfile_N59) );
  MUX2_X2 U14417 ( .A(decode_regfile_fpregs_30__1_), .B(
        decode_regfile_fpregs_31__1_), .S(n10824), .Z(n9816) );
  MUX2_X2 U14418 ( .A(decode_regfile_fpregs_28__1_), .B(
        decode_regfile_fpregs_29__1_), .S(n10825), .Z(n9817) );
  MUX2_X2 U14419 ( .A(n9817), .B(n9816), .S(n10903), .Z(n9818) );
  MUX2_X2 U14420 ( .A(decode_regfile_fpregs_26__1_), .B(
        decode_regfile_fpregs_27__1_), .S(n10825), .Z(n9819) );
  MUX2_X2 U14421 ( .A(decode_regfile_fpregs_24__1_), .B(
        decode_regfile_fpregs_25__1_), .S(n10825), .Z(n9820) );
  MUX2_X2 U14422 ( .A(n9820), .B(n9819), .S(n10903), .Z(n9821) );
  MUX2_X2 U14423 ( .A(n9821), .B(n9818), .S(n10933), .Z(n9822) );
  MUX2_X2 U14424 ( .A(decode_regfile_fpregs_22__1_), .B(
        decode_regfile_fpregs_23__1_), .S(n10825), .Z(n9823) );
  MUX2_X2 U14425 ( .A(decode_regfile_fpregs_20__1_), .B(
        decode_regfile_fpregs_21__1_), .S(n10825), .Z(n9824) );
  MUX2_X2 U14426 ( .A(n9824), .B(n9823), .S(n10903), .Z(n9825) );
  MUX2_X2 U14427 ( .A(decode_regfile_fpregs_18__1_), .B(
        decode_regfile_fpregs_19__1_), .S(n10825), .Z(n9826) );
  MUX2_X2 U14428 ( .A(decode_regfile_fpregs_16__1_), .B(
        decode_regfile_fpregs_17__1_), .S(n10825), .Z(n9827) );
  MUX2_X2 U14429 ( .A(n9827), .B(n9826), .S(n10903), .Z(n9828) );
  MUX2_X2 U14430 ( .A(n9828), .B(n9825), .S(n10933), .Z(n9829) );
  MUX2_X2 U14431 ( .A(n9829), .B(n9822), .S(n10949), .Z(n9830) );
  MUX2_X2 U14432 ( .A(decode_regfile_fpregs_14__1_), .B(
        decode_regfile_fpregs_15__1_), .S(n10825), .Z(n9831) );
  MUX2_X2 U14433 ( .A(decode_regfile_fpregs_12__1_), .B(
        decode_regfile_fpregs_13__1_), .S(n10825), .Z(n9832) );
  MUX2_X2 U14434 ( .A(n9832), .B(n9831), .S(n10903), .Z(n9833) );
  MUX2_X2 U14435 ( .A(decode_regfile_fpregs_10__1_), .B(
        decode_regfile_fpregs_11__1_), .S(n10825), .Z(n9834) );
  MUX2_X2 U14436 ( .A(decode_regfile_fpregs_8__1_), .B(
        decode_regfile_fpregs_9__1_), .S(n10825), .Z(n9835) );
  MUX2_X2 U14437 ( .A(n9835), .B(n9834), .S(n10903), .Z(n9836) );
  MUX2_X2 U14438 ( .A(n9836), .B(n9833), .S(n10933), .Z(n9837) );
  MUX2_X2 U14439 ( .A(decode_regfile_fpregs_6__1_), .B(
        decode_regfile_fpregs_7__1_), .S(n10826), .Z(n9838) );
  MUX2_X2 U14440 ( .A(decode_regfile_fpregs_4__1_), .B(
        decode_regfile_fpregs_5__1_), .S(n10826), .Z(n9839) );
  MUX2_X2 U14441 ( .A(n9839), .B(n9838), .S(n10904), .Z(n9840) );
  MUX2_X2 U14442 ( .A(decode_regfile_fpregs_2__1_), .B(
        decode_regfile_fpregs_3__1_), .S(n10826), .Z(n9841) );
  MUX2_X2 U14443 ( .A(decode_regfile_fpregs_0__1_), .B(
        decode_regfile_fpregs_1__1_), .S(n10826), .Z(n9842) );
  MUX2_X2 U14444 ( .A(n9842), .B(n9841), .S(n10904), .Z(n9843) );
  MUX2_X2 U14445 ( .A(n9843), .B(n9840), .S(n10934), .Z(n9844) );
  MUX2_X2 U14446 ( .A(n9844), .B(n9837), .S(n10949), .Z(n9845) );
  MUX2_X2 U14447 ( .A(n9845), .B(n9830), .S(n10958), .Z(decode_regfile_N58) );
  MUX2_X2 U14448 ( .A(decode_regfile_fpregs_30__2_), .B(
        decode_regfile_fpregs_31__2_), .S(n10826), .Z(n9846) );
  MUX2_X2 U14449 ( .A(decode_regfile_fpregs_28__2_), .B(
        decode_regfile_fpregs_29__2_), .S(n10826), .Z(n9847) );
  MUX2_X2 U14450 ( .A(n9847), .B(n9846), .S(n10904), .Z(n9848) );
  MUX2_X2 U14451 ( .A(decode_regfile_fpregs_26__2_), .B(
        decode_regfile_fpregs_27__2_), .S(n10826), .Z(n9849) );
  MUX2_X2 U14452 ( .A(decode_regfile_fpregs_24__2_), .B(
        decode_regfile_fpregs_25__2_), .S(n10826), .Z(n9850) );
  MUX2_X2 U14453 ( .A(n9850), .B(n9849), .S(n10904), .Z(n9851) );
  MUX2_X2 U14454 ( .A(n9851), .B(n9848), .S(n10934), .Z(n9852) );
  MUX2_X2 U14455 ( .A(decode_regfile_fpregs_22__2_), .B(
        decode_regfile_fpregs_23__2_), .S(n10826), .Z(n9853) );
  MUX2_X2 U14456 ( .A(decode_regfile_fpregs_20__2_), .B(
        decode_regfile_fpregs_21__2_), .S(n10826), .Z(n9854) );
  MUX2_X2 U14457 ( .A(n9854), .B(n9853), .S(n10904), .Z(n9855) );
  MUX2_X2 U14458 ( .A(decode_regfile_fpregs_18__2_), .B(
        decode_regfile_fpregs_19__2_), .S(n10826), .Z(n9856) );
  MUX2_X2 U14459 ( .A(decode_regfile_fpregs_16__2_), .B(
        decode_regfile_fpregs_17__2_), .S(n10827), .Z(n9857) );
  MUX2_X2 U14460 ( .A(n9857), .B(n9856), .S(n10904), .Z(n9858) );
  MUX2_X2 U14461 ( .A(n9858), .B(n9855), .S(n10934), .Z(n9859) );
  MUX2_X2 U14462 ( .A(n9859), .B(n9852), .S(n10949), .Z(n9860) );
  MUX2_X2 U14463 ( .A(decode_regfile_fpregs_14__2_), .B(
        decode_regfile_fpregs_15__2_), .S(n10827), .Z(n9861) );
  MUX2_X2 U14464 ( .A(decode_regfile_fpregs_12__2_), .B(
        decode_regfile_fpregs_13__2_), .S(n10827), .Z(n9862) );
  MUX2_X2 U14465 ( .A(n9862), .B(n9861), .S(n10904), .Z(n9863) );
  MUX2_X2 U14466 ( .A(decode_regfile_fpregs_10__2_), .B(
        decode_regfile_fpregs_11__2_), .S(n10827), .Z(n9864) );
  MUX2_X2 U14467 ( .A(decode_regfile_fpregs_8__2_), .B(
        decode_regfile_fpregs_9__2_), .S(n10827), .Z(n9865) );
  MUX2_X2 U14468 ( .A(n9865), .B(n9864), .S(n10904), .Z(n9866) );
  MUX2_X2 U14469 ( .A(n9866), .B(n9863), .S(n10934), .Z(n9867) );
  MUX2_X2 U14470 ( .A(decode_regfile_fpregs_6__2_), .B(
        decode_regfile_fpregs_7__2_), .S(n10827), .Z(n9868) );
  MUX2_X2 U14471 ( .A(decode_regfile_fpregs_4__2_), .B(
        decode_regfile_fpregs_5__2_), .S(n10827), .Z(n9869) );
  MUX2_X2 U14472 ( .A(n9869), .B(n9868), .S(n10904), .Z(n9870) );
  MUX2_X2 U14473 ( .A(decode_regfile_fpregs_2__2_), .B(
        decode_regfile_fpregs_3__2_), .S(n10827), .Z(n9871) );
  MUX2_X2 U14474 ( .A(decode_regfile_fpregs_0__2_), .B(
        decode_regfile_fpregs_1__2_), .S(n10827), .Z(n9872) );
  MUX2_X2 U14475 ( .A(n9872), .B(n9871), .S(n10904), .Z(n9873) );
  MUX2_X2 U14476 ( .A(n9873), .B(n9870), .S(n10934), .Z(n9874) );
  MUX2_X2 U14477 ( .A(n9874), .B(n9867), .S(n10949), .Z(n9875) );
  MUX2_X2 U14478 ( .A(n9875), .B(n9860), .S(n10958), .Z(decode_regfile_N57) );
  MUX2_X2 U14479 ( .A(decode_regfile_fpregs_30__3_), .B(
        decode_regfile_fpregs_31__3_), .S(n10827), .Z(n9876) );
  MUX2_X2 U14480 ( .A(decode_regfile_fpregs_28__3_), .B(
        decode_regfile_fpregs_29__3_), .S(n10827), .Z(n9877) );
  MUX2_X2 U14481 ( .A(n9877), .B(n9876), .S(n10904), .Z(n9878) );
  MUX2_X2 U14482 ( .A(decode_regfile_fpregs_26__3_), .B(
        decode_regfile_fpregs_27__3_), .S(n10828), .Z(n9879) );
  MUX2_X2 U14483 ( .A(decode_regfile_fpregs_24__3_), .B(
        decode_regfile_fpregs_25__3_), .S(n10828), .Z(n9880) );
  MUX2_X2 U14484 ( .A(n9880), .B(n9879), .S(n10905), .Z(n9881) );
  MUX2_X2 U14485 ( .A(n9881), .B(n9878), .S(n10934), .Z(n9882) );
  MUX2_X2 U14486 ( .A(decode_regfile_fpregs_22__3_), .B(
        decode_regfile_fpregs_23__3_), .S(n10828), .Z(n9883) );
  MUX2_X2 U14487 ( .A(decode_regfile_fpregs_20__3_), .B(
        decode_regfile_fpregs_21__3_), .S(n10828), .Z(n9884) );
  MUX2_X2 U14488 ( .A(n9884), .B(n9883), .S(n10905), .Z(n9885) );
  MUX2_X2 U14489 ( .A(decode_regfile_fpregs_18__3_), .B(
        decode_regfile_fpregs_19__3_), .S(n10828), .Z(n9886) );
  MUX2_X2 U14490 ( .A(decode_regfile_fpregs_16__3_), .B(
        decode_regfile_fpregs_17__3_), .S(n10828), .Z(n9887) );
  MUX2_X2 U14491 ( .A(n9887), .B(n9886), .S(n10905), .Z(n9888) );
  MUX2_X2 U14492 ( .A(n9888), .B(n9885), .S(n10934), .Z(n9889) );
  MUX2_X2 U14493 ( .A(n9889), .B(n9882), .S(n10949), .Z(n9890) );
  MUX2_X2 U14494 ( .A(decode_regfile_fpregs_14__3_), .B(
        decode_regfile_fpregs_15__3_), .S(n10828), .Z(n9891) );
  MUX2_X2 U14495 ( .A(decode_regfile_fpregs_12__3_), .B(
        decode_regfile_fpregs_13__3_), .S(n10828), .Z(n9892) );
  MUX2_X2 U14496 ( .A(n9892), .B(n9891), .S(n10905), .Z(n9893) );
  MUX2_X2 U14497 ( .A(decode_regfile_fpregs_10__3_), .B(
        decode_regfile_fpregs_11__3_), .S(n10828), .Z(n9894) );
  MUX2_X2 U14498 ( .A(decode_regfile_fpregs_8__3_), .B(
        decode_regfile_fpregs_9__3_), .S(n10828), .Z(n9895) );
  MUX2_X2 U14499 ( .A(n9895), .B(n9894), .S(n10905), .Z(n9896) );
  MUX2_X2 U14500 ( .A(n9896), .B(n9893), .S(n10934), .Z(n9897) );
  MUX2_X2 U14501 ( .A(decode_regfile_fpregs_6__3_), .B(
        decode_regfile_fpregs_7__3_), .S(n10828), .Z(n9898) );
  MUX2_X2 U14502 ( .A(decode_regfile_fpregs_4__3_), .B(
        decode_regfile_fpregs_5__3_), .S(n10829), .Z(n9899) );
  MUX2_X2 U14503 ( .A(n9899), .B(n9898), .S(n10905), .Z(n9900) );
  MUX2_X2 U14504 ( .A(decode_regfile_fpregs_2__3_), .B(
        decode_regfile_fpregs_3__3_), .S(n10829), .Z(n9901) );
  MUX2_X2 U14505 ( .A(decode_regfile_fpregs_0__3_), .B(
        decode_regfile_fpregs_1__3_), .S(n10829), .Z(n9902) );
  MUX2_X2 U14506 ( .A(n9902), .B(n9901), .S(n10905), .Z(n9903) );
  MUX2_X2 U14507 ( .A(n9903), .B(n9900), .S(n10934), .Z(n9904) );
  MUX2_X2 U14508 ( .A(n9904), .B(n9897), .S(n10949), .Z(n9905) );
  MUX2_X2 U14509 ( .A(n9905), .B(n9890), .S(n10958), .Z(decode_regfile_N56) );
  MUX2_X2 U14510 ( .A(decode_regfile_fpregs_30__4_), .B(
        decode_regfile_fpregs_31__4_), .S(n10829), .Z(n9906) );
  MUX2_X2 U14511 ( .A(decode_regfile_fpregs_28__4_), .B(
        decode_regfile_fpregs_29__4_), .S(n10829), .Z(n9907) );
  MUX2_X2 U14512 ( .A(n9907), .B(n9906), .S(n10905), .Z(n9908) );
  MUX2_X2 U14513 ( .A(decode_regfile_fpregs_26__4_), .B(
        decode_regfile_fpregs_27__4_), .S(n10829), .Z(n9909) );
  MUX2_X2 U14514 ( .A(decode_regfile_fpregs_24__4_), .B(
        decode_regfile_fpregs_25__4_), .S(n10829), .Z(n9910) );
  MUX2_X2 U14515 ( .A(n9910), .B(n9909), .S(n10905), .Z(n9911) );
  MUX2_X2 U14516 ( .A(n9911), .B(n9908), .S(n10934), .Z(n9912) );
  MUX2_X2 U14517 ( .A(decode_regfile_fpregs_22__4_), .B(
        decode_regfile_fpregs_23__4_), .S(n10829), .Z(n9913) );
  MUX2_X2 U14518 ( .A(decode_regfile_fpregs_20__4_), .B(
        decode_regfile_fpregs_21__4_), .S(n10829), .Z(n9914) );
  MUX2_X2 U14519 ( .A(n9914), .B(n9913), .S(n10905), .Z(n9915) );
  MUX2_X2 U14520 ( .A(decode_regfile_fpregs_18__4_), .B(
        decode_regfile_fpregs_19__4_), .S(n10829), .Z(n9916) );
  MUX2_X2 U14521 ( .A(decode_regfile_fpregs_16__4_), .B(
        decode_regfile_fpregs_17__4_), .S(n10829), .Z(n9917) );
  MUX2_X2 U14522 ( .A(n9917), .B(n9916), .S(n10905), .Z(n9918) );
  MUX2_X2 U14523 ( .A(n9918), .B(n9915), .S(n10934), .Z(n9919) );
  MUX2_X2 U14524 ( .A(n9919), .B(n9912), .S(n10949), .Z(n9920) );
  MUX2_X2 U14525 ( .A(decode_regfile_fpregs_14__4_), .B(
        decode_regfile_fpregs_15__4_), .S(n10830), .Z(n9921) );
  MUX2_X2 U14526 ( .A(decode_regfile_fpregs_12__4_), .B(
        decode_regfile_fpregs_13__4_), .S(n10830), .Z(n9922) );
  MUX2_X2 U14527 ( .A(n9922), .B(n9921), .S(n10906), .Z(n9923) );
  MUX2_X2 U14528 ( .A(decode_regfile_fpregs_10__4_), .B(
        decode_regfile_fpregs_11__4_), .S(n10830), .Z(n9924) );
  MUX2_X2 U14529 ( .A(decode_regfile_fpregs_8__4_), .B(
        decode_regfile_fpregs_9__4_), .S(n10830), .Z(n9925) );
  MUX2_X2 U14530 ( .A(n9925), .B(n9924), .S(n10906), .Z(n9926) );
  MUX2_X2 U14531 ( .A(n9926), .B(n9923), .S(n10935), .Z(n9927) );
  MUX2_X2 U14532 ( .A(decode_regfile_fpregs_6__4_), .B(
        decode_regfile_fpregs_7__4_), .S(n10830), .Z(n9928) );
  MUX2_X2 U14533 ( .A(decode_regfile_fpregs_4__4_), .B(
        decode_regfile_fpregs_5__4_), .S(n10830), .Z(n9929) );
  MUX2_X2 U14534 ( .A(n9929), .B(n9928), .S(n10906), .Z(n9930) );
  MUX2_X2 U14535 ( .A(decode_regfile_fpregs_2__4_), .B(
        decode_regfile_fpregs_3__4_), .S(n10830), .Z(n9931) );
  MUX2_X2 U14536 ( .A(decode_regfile_fpregs_0__4_), .B(
        decode_regfile_fpregs_1__4_), .S(n10830), .Z(n9932) );
  MUX2_X2 U14537 ( .A(n9932), .B(n9931), .S(n10906), .Z(n9933) );
  MUX2_X2 U14538 ( .A(n9933), .B(n9930), .S(n10935), .Z(n9934) );
  MUX2_X2 U14539 ( .A(n9934), .B(n9927), .S(n10950), .Z(n9935) );
  MUX2_X2 U14540 ( .A(n9935), .B(n9920), .S(n10958), .Z(decode_regfile_N55) );
  MUX2_X2 U14541 ( .A(decode_regfile_fpregs_30__5_), .B(
        decode_regfile_fpregs_31__5_), .S(n10830), .Z(n9936) );
  MUX2_X2 U14542 ( .A(decode_regfile_fpregs_28__5_), .B(
        decode_regfile_fpregs_29__5_), .S(n10830), .Z(n9937) );
  MUX2_X2 U14543 ( .A(n9937), .B(n9936), .S(n10906), .Z(n9938) );
  MUX2_X2 U14544 ( .A(decode_regfile_fpregs_26__5_), .B(
        decode_regfile_fpregs_27__5_), .S(n10830), .Z(n9939) );
  MUX2_X2 U14545 ( .A(decode_regfile_fpregs_24__5_), .B(
        decode_regfile_fpregs_25__5_), .S(n10831), .Z(n9940) );
  MUX2_X2 U14546 ( .A(n9940), .B(n9939), .S(n10906), .Z(n9941) );
  MUX2_X2 U14547 ( .A(n9941), .B(n9938), .S(n10935), .Z(n9942) );
  MUX2_X2 U14548 ( .A(decode_regfile_fpregs_22__5_), .B(
        decode_regfile_fpregs_23__5_), .S(n10831), .Z(n9943) );
  MUX2_X2 U14549 ( .A(decode_regfile_fpregs_20__5_), .B(
        decode_regfile_fpregs_21__5_), .S(n10831), .Z(n9944) );
  MUX2_X2 U14550 ( .A(n9944), .B(n9943), .S(n10906), .Z(n9945) );
  MUX2_X2 U14551 ( .A(decode_regfile_fpregs_18__5_), .B(
        decode_regfile_fpregs_19__5_), .S(n10831), .Z(n9946) );
  MUX2_X2 U14552 ( .A(decode_regfile_fpregs_16__5_), .B(
        decode_regfile_fpregs_17__5_), .S(n10831), .Z(n9947) );
  MUX2_X2 U14553 ( .A(n9947), .B(n9946), .S(n10906), .Z(n9948) );
  MUX2_X2 U14554 ( .A(n9948), .B(n9945), .S(n10935), .Z(n9949) );
  MUX2_X2 U14555 ( .A(n9949), .B(n9942), .S(n10950), .Z(n9950) );
  MUX2_X2 U14556 ( .A(decode_regfile_fpregs_14__5_), .B(
        decode_regfile_fpregs_15__5_), .S(n10831), .Z(n9951) );
  MUX2_X2 U14557 ( .A(decode_regfile_fpregs_12__5_), .B(
        decode_regfile_fpregs_13__5_), .S(n10831), .Z(n9952) );
  MUX2_X2 U14558 ( .A(n9952), .B(n9951), .S(n10906), .Z(n9953) );
  MUX2_X2 U14559 ( .A(decode_regfile_fpregs_10__5_), .B(
        decode_regfile_fpregs_11__5_), .S(n10831), .Z(n9954) );
  MUX2_X2 U14560 ( .A(decode_regfile_fpregs_8__5_), .B(
        decode_regfile_fpregs_9__5_), .S(n10831), .Z(n9955) );
  MUX2_X2 U14561 ( .A(n9955), .B(n9954), .S(n10906), .Z(n9956) );
  MUX2_X2 U14562 ( .A(n9956), .B(n9953), .S(n10935), .Z(n9957) );
  MUX2_X2 U14563 ( .A(decode_regfile_fpregs_6__5_), .B(
        decode_regfile_fpregs_7__5_), .S(n10831), .Z(n9958) );
  MUX2_X2 U14564 ( .A(decode_regfile_fpregs_4__5_), .B(
        decode_regfile_fpregs_5__5_), .S(n10831), .Z(n9959) );
  MUX2_X2 U14565 ( .A(n9959), .B(n9958), .S(n10906), .Z(n9960) );
  MUX2_X2 U14566 ( .A(decode_regfile_fpregs_2__5_), .B(
        decode_regfile_fpregs_3__5_), .S(n10832), .Z(n9961) );
  MUX2_X2 U14567 ( .A(decode_regfile_fpregs_0__5_), .B(
        decode_regfile_fpregs_1__5_), .S(n10832), .Z(n9962) );
  MUX2_X2 U14568 ( .A(n9962), .B(n9961), .S(n10907), .Z(n9963) );
  MUX2_X2 U14569 ( .A(n9963), .B(n9960), .S(n10935), .Z(n9964) );
  MUX2_X2 U14570 ( .A(n9964), .B(n9957), .S(n10950), .Z(n9965) );
  MUX2_X2 U14571 ( .A(n9965), .B(n9950), .S(n10958), .Z(decode_regfile_N54) );
  MUX2_X2 U14572 ( .A(decode_regfile_fpregs_30__6_), .B(
        decode_regfile_fpregs_31__6_), .S(n10832), .Z(n9966) );
  MUX2_X2 U14573 ( .A(decode_regfile_fpregs_28__6_), .B(
        decode_regfile_fpregs_29__6_), .S(n10832), .Z(n9967) );
  MUX2_X2 U14574 ( .A(n9967), .B(n9966), .S(n10907), .Z(n9968) );
  MUX2_X2 U14575 ( .A(decode_regfile_fpregs_26__6_), .B(
        decode_regfile_fpregs_27__6_), .S(n10832), .Z(n9969) );
  MUX2_X2 U14576 ( .A(decode_regfile_fpregs_24__6_), .B(
        decode_regfile_fpregs_25__6_), .S(n10832), .Z(n9970) );
  MUX2_X2 U14577 ( .A(n9970), .B(n9969), .S(n10907), .Z(n9971) );
  MUX2_X2 U14578 ( .A(n9971), .B(n9968), .S(n10935), .Z(n9972) );
  MUX2_X2 U14579 ( .A(decode_regfile_fpregs_22__6_), .B(
        decode_regfile_fpregs_23__6_), .S(n10832), .Z(n9973) );
  MUX2_X2 U14580 ( .A(decode_regfile_fpregs_20__6_), .B(
        decode_regfile_fpregs_21__6_), .S(n10832), .Z(n9974) );
  MUX2_X2 U14581 ( .A(n9974), .B(n9973), .S(n10907), .Z(n9975) );
  MUX2_X2 U14582 ( .A(decode_regfile_fpregs_18__6_), .B(
        decode_regfile_fpregs_19__6_), .S(n10832), .Z(n9976) );
  MUX2_X2 U14583 ( .A(decode_regfile_fpregs_16__6_), .B(
        decode_regfile_fpregs_17__6_), .S(n10832), .Z(n9977) );
  MUX2_X2 U14584 ( .A(n9977), .B(n9976), .S(n10907), .Z(n9978) );
  MUX2_X2 U14585 ( .A(n9978), .B(n9975), .S(n10935), .Z(n9979) );
  MUX2_X2 U14586 ( .A(n9979), .B(n9972), .S(n10950), .Z(n9980) );
  MUX2_X2 U14587 ( .A(decode_regfile_fpregs_14__6_), .B(
        decode_regfile_fpregs_15__6_), .S(n10832), .Z(n9981) );
  MUX2_X2 U14588 ( .A(decode_regfile_fpregs_12__6_), .B(
        decode_regfile_fpregs_13__6_), .S(n10833), .Z(n9982) );
  MUX2_X2 U14589 ( .A(n9982), .B(n9981), .S(n10907), .Z(n9983) );
  MUX2_X2 U14590 ( .A(decode_regfile_fpregs_10__6_), .B(
        decode_regfile_fpregs_11__6_), .S(n10833), .Z(n9984) );
  MUX2_X2 U14591 ( .A(decode_regfile_fpregs_8__6_), .B(
        decode_regfile_fpregs_9__6_), .S(n10833), .Z(n9985) );
  MUX2_X2 U14592 ( .A(n9985), .B(n9984), .S(n10907), .Z(n9986) );
  MUX2_X2 U14593 ( .A(n9986), .B(n9983), .S(n10935), .Z(n9987) );
  MUX2_X2 U14594 ( .A(decode_regfile_fpregs_6__6_), .B(
        decode_regfile_fpregs_7__6_), .S(n10833), .Z(n9988) );
  MUX2_X2 U14595 ( .A(decode_regfile_fpregs_4__6_), .B(
        decode_regfile_fpregs_5__6_), .S(n10833), .Z(n9989) );
  MUX2_X2 U14596 ( .A(n9989), .B(n9988), .S(n10907), .Z(n9990) );
  MUX2_X2 U14597 ( .A(decode_regfile_fpregs_2__6_), .B(
        decode_regfile_fpregs_3__6_), .S(n10833), .Z(n9991) );
  MUX2_X2 U14598 ( .A(decode_regfile_fpregs_0__6_), .B(
        decode_regfile_fpregs_1__6_), .S(n10833), .Z(n9992) );
  MUX2_X2 U14599 ( .A(n9992), .B(n9991), .S(n10907), .Z(n9993) );
  MUX2_X2 U14600 ( .A(n9993), .B(n9990), .S(n10935), .Z(n9994) );
  MUX2_X2 U14601 ( .A(n9994), .B(n9987), .S(n10950), .Z(n9995) );
  MUX2_X2 U14602 ( .A(n9995), .B(n9980), .S(n10958), .Z(decode_regfile_N53) );
  MUX2_X2 U14603 ( .A(decode_regfile_fpregs_30__7_), .B(
        decode_regfile_fpregs_31__7_), .S(n10833), .Z(n9996) );
  MUX2_X2 U14604 ( .A(decode_regfile_fpregs_28__7_), .B(
        decode_regfile_fpregs_29__7_), .S(n10833), .Z(n9997) );
  MUX2_X2 U14605 ( .A(n9997), .B(n9996), .S(n10907), .Z(n9998) );
  MUX2_X2 U14606 ( .A(decode_regfile_fpregs_26__7_), .B(
        decode_regfile_fpregs_27__7_), .S(n10833), .Z(n9999) );
  MUX2_X2 U14607 ( .A(decode_regfile_fpregs_24__7_), .B(
        decode_regfile_fpregs_25__7_), .S(n10833), .Z(n10000) );
  MUX2_X2 U14608 ( .A(n10000), .B(n9999), .S(n10907), .Z(n10001) );
  MUX2_X2 U14609 ( .A(n10001), .B(n9998), .S(n10935), .Z(n10002) );
  MUX2_X2 U14610 ( .A(decode_regfile_fpregs_22__7_), .B(
        decode_regfile_fpregs_23__7_), .S(n10834), .Z(n10003) );
  MUX2_X2 U14611 ( .A(decode_regfile_fpregs_20__7_), .B(
        decode_regfile_fpregs_21__7_), .S(n10834), .Z(n10004) );
  MUX2_X2 U14612 ( .A(n10004), .B(n10003), .S(n10908), .Z(n10005) );
  MUX2_X2 U14613 ( .A(decode_regfile_fpregs_18__7_), .B(
        decode_regfile_fpregs_19__7_), .S(n10834), .Z(n10006) );
  MUX2_X2 U14614 ( .A(decode_regfile_fpregs_16__7_), .B(
        decode_regfile_fpregs_17__7_), .S(n10834), .Z(n10007) );
  MUX2_X2 U14615 ( .A(n10007), .B(n10006), .S(n10908), .Z(n10008) );
  MUX2_X2 U14616 ( .A(n10008), .B(n10005), .S(n10936), .Z(n10009) );
  MUX2_X2 U14617 ( .A(n10009), .B(n10002), .S(n10950), .Z(n10010) );
  MUX2_X2 U14618 ( .A(decode_regfile_fpregs_14__7_), .B(
        decode_regfile_fpregs_15__7_), .S(n10834), .Z(n10011) );
  MUX2_X2 U14619 ( .A(decode_regfile_fpregs_12__7_), .B(
        decode_regfile_fpregs_13__7_), .S(n10834), .Z(n10012) );
  MUX2_X2 U14620 ( .A(n10012), .B(n10011), .S(n10908), .Z(n10013) );
  MUX2_X2 U14621 ( .A(decode_regfile_fpregs_10__7_), .B(
        decode_regfile_fpregs_11__7_), .S(n10834), .Z(n10014) );
  MUX2_X2 U14622 ( .A(decode_regfile_fpregs_8__7_), .B(
        decode_regfile_fpregs_9__7_), .S(n10834), .Z(n10015) );
  MUX2_X2 U14623 ( .A(n10015), .B(n10014), .S(n10908), .Z(n10016) );
  MUX2_X2 U14624 ( .A(n10016), .B(n10013), .S(n10936), .Z(n10017) );
  MUX2_X2 U14625 ( .A(decode_regfile_fpregs_6__7_), .B(
        decode_regfile_fpregs_7__7_), .S(n10834), .Z(n10018) );
  MUX2_X2 U14626 ( .A(decode_regfile_fpregs_4__7_), .B(
        decode_regfile_fpregs_5__7_), .S(n10834), .Z(n10019) );
  MUX2_X2 U14627 ( .A(n10019), .B(n10018), .S(n10908), .Z(n10020) );
  MUX2_X2 U14628 ( .A(decode_regfile_fpregs_2__7_), .B(
        decode_regfile_fpregs_3__7_), .S(n10834), .Z(n10021) );
  MUX2_X2 U14629 ( .A(decode_regfile_fpregs_0__7_), .B(
        decode_regfile_fpregs_1__7_), .S(n10835), .Z(n10022) );
  MUX2_X2 U14630 ( .A(n10022), .B(n10021), .S(n10908), .Z(n10023) );
  MUX2_X2 U14631 ( .A(n10023), .B(n10020), .S(n10936), .Z(n10024) );
  MUX2_X2 U14632 ( .A(n10024), .B(n10017), .S(n10950), .Z(n10025) );
  MUX2_X2 U14633 ( .A(n10025), .B(n10010), .S(n10958), .Z(decode_regfile_N52)
         );
  MUX2_X2 U14634 ( .A(decode_regfile_fpregs_30__8_), .B(
        decode_regfile_fpregs_31__8_), .S(n10835), .Z(n10026) );
  MUX2_X2 U14635 ( .A(decode_regfile_fpregs_28__8_), .B(
        decode_regfile_fpregs_29__8_), .S(n10835), .Z(n10027) );
  MUX2_X2 U14636 ( .A(n10027), .B(n10026), .S(n10908), .Z(n10028) );
  MUX2_X2 U14637 ( .A(decode_regfile_fpregs_26__8_), .B(
        decode_regfile_fpregs_27__8_), .S(n10835), .Z(n10029) );
  MUX2_X2 U14638 ( .A(decode_regfile_fpregs_24__8_), .B(
        decode_regfile_fpregs_25__8_), .S(n10835), .Z(n10030) );
  MUX2_X2 U14639 ( .A(n10030), .B(n10029), .S(n10908), .Z(n10031) );
  MUX2_X2 U14640 ( .A(n10031), .B(n10028), .S(n10936), .Z(n10032) );
  MUX2_X2 U14641 ( .A(decode_regfile_fpregs_22__8_), .B(
        decode_regfile_fpregs_23__8_), .S(n10835), .Z(n10033) );
  MUX2_X2 U14642 ( .A(decode_regfile_fpregs_20__8_), .B(
        decode_regfile_fpregs_21__8_), .S(n10835), .Z(n10034) );
  MUX2_X2 U14643 ( .A(n10034), .B(n10033), .S(n10908), .Z(n10035) );
  MUX2_X2 U14644 ( .A(decode_regfile_fpregs_18__8_), .B(
        decode_regfile_fpregs_19__8_), .S(n10835), .Z(n10036) );
  MUX2_X2 U14645 ( .A(decode_regfile_fpregs_16__8_), .B(
        decode_regfile_fpregs_17__8_), .S(n10835), .Z(n10037) );
  MUX2_X2 U14646 ( .A(n10037), .B(n10036), .S(n10908), .Z(n10038) );
  MUX2_X2 U14647 ( .A(n10038), .B(n10035), .S(n10936), .Z(n10039) );
  MUX2_X2 U14648 ( .A(n10039), .B(n10032), .S(n10950), .Z(n10040) );
  MUX2_X2 U14649 ( .A(decode_regfile_fpregs_14__8_), .B(
        decode_regfile_fpregs_15__8_), .S(n10835), .Z(n10041) );
  MUX2_X2 U14650 ( .A(decode_regfile_fpregs_12__8_), .B(
        decode_regfile_fpregs_13__8_), .S(n10835), .Z(n10042) );
  MUX2_X2 U14651 ( .A(n10042), .B(n10041), .S(n10908), .Z(n10043) );
  MUX2_X2 U14652 ( .A(decode_regfile_fpregs_10__8_), .B(
        decode_regfile_fpregs_11__8_), .S(n10836), .Z(n10044) );
  MUX2_X2 U14653 ( .A(decode_regfile_fpregs_8__8_), .B(
        decode_regfile_fpregs_9__8_), .S(n10836), .Z(n10045) );
  MUX2_X2 U14654 ( .A(n10045), .B(n10044), .S(n10909), .Z(n10046) );
  MUX2_X2 U14655 ( .A(n10046), .B(n10043), .S(n10936), .Z(n10047) );
  MUX2_X2 U14656 ( .A(decode_regfile_fpregs_6__8_), .B(
        decode_regfile_fpregs_7__8_), .S(n10836), .Z(n10048) );
  MUX2_X2 U14657 ( .A(decode_regfile_fpregs_4__8_), .B(
        decode_regfile_fpregs_5__8_), .S(n10836), .Z(n10049) );
  MUX2_X2 U14658 ( .A(n10049), .B(n10048), .S(n10909), .Z(n10050) );
  MUX2_X2 U14659 ( .A(decode_regfile_fpregs_2__8_), .B(
        decode_regfile_fpregs_3__8_), .S(n10836), .Z(n10051) );
  MUX2_X2 U14660 ( .A(decode_regfile_fpregs_0__8_), .B(
        decode_regfile_fpregs_1__8_), .S(n10836), .Z(n10052) );
  MUX2_X2 U14661 ( .A(n10052), .B(n10051), .S(n10909), .Z(n10053) );
  MUX2_X2 U14662 ( .A(n10053), .B(n10050), .S(n10936), .Z(n10054) );
  MUX2_X2 U14663 ( .A(n10054), .B(n10047), .S(n10950), .Z(n10055) );
  MUX2_X2 U14664 ( .A(n10055), .B(n10040), .S(n10958), .Z(decode_regfile_N51)
         );
  MUX2_X2 U14665 ( .A(decode_regfile_fpregs_30__9_), .B(
        decode_regfile_fpregs_31__9_), .S(n10836), .Z(n10056) );
  MUX2_X2 U14666 ( .A(decode_regfile_fpregs_28__9_), .B(
        decode_regfile_fpregs_29__9_), .S(n10836), .Z(n10057) );
  MUX2_X2 U14667 ( .A(n10057), .B(n10056), .S(n10909), .Z(n10058) );
  MUX2_X2 U14668 ( .A(decode_regfile_fpregs_26__9_), .B(
        decode_regfile_fpregs_27__9_), .S(n10836), .Z(n10059) );
  MUX2_X2 U14669 ( .A(decode_regfile_fpregs_24__9_), .B(
        decode_regfile_fpregs_25__9_), .S(n10836), .Z(n10060) );
  MUX2_X2 U14670 ( .A(n10060), .B(n10059), .S(n10909), .Z(n10061) );
  MUX2_X2 U14671 ( .A(n10061), .B(n10058), .S(n10936), .Z(n10062) );
  MUX2_X2 U14672 ( .A(decode_regfile_fpregs_22__9_), .B(
        decode_regfile_fpregs_23__9_), .S(n10836), .Z(n10063) );
  MUX2_X2 U14673 ( .A(decode_regfile_fpregs_20__9_), .B(
        decode_regfile_fpregs_21__9_), .S(n10837), .Z(n10064) );
  MUX2_X2 U14674 ( .A(n10064), .B(n10063), .S(n10909), .Z(n10065) );
  MUX2_X2 U14675 ( .A(decode_regfile_fpregs_18__9_), .B(
        decode_regfile_fpregs_19__9_), .S(n10837), .Z(n10066) );
  MUX2_X2 U14676 ( .A(decode_regfile_fpregs_16__9_), .B(
        decode_regfile_fpregs_17__9_), .S(n10837), .Z(n10067) );
  MUX2_X2 U14677 ( .A(n10067), .B(n10066), .S(n10909), .Z(n10068) );
  MUX2_X2 U14678 ( .A(n10068), .B(n10065), .S(n10936), .Z(n10069) );
  MUX2_X2 U14679 ( .A(n10069), .B(n10062), .S(n10950), .Z(n10070) );
  MUX2_X2 U14680 ( .A(decode_regfile_fpregs_14__9_), .B(
        decode_regfile_fpregs_15__9_), .S(n10837), .Z(n10071) );
  MUX2_X2 U14681 ( .A(decode_regfile_fpregs_12__9_), .B(
        decode_regfile_fpregs_13__9_), .S(n10837), .Z(n10072) );
  MUX2_X2 U14682 ( .A(n10072), .B(n10071), .S(n10909), .Z(n10073) );
  MUX2_X2 U14683 ( .A(decode_regfile_fpregs_10__9_), .B(
        decode_regfile_fpregs_11__9_), .S(n10837), .Z(n10074) );
  MUX2_X2 U14684 ( .A(decode_regfile_fpregs_8__9_), .B(
        decode_regfile_fpregs_9__9_), .S(n10837), .Z(n10075) );
  MUX2_X2 U14685 ( .A(n10075), .B(n10074), .S(n10909), .Z(n10076) );
  MUX2_X2 U14686 ( .A(n10076), .B(n10073), .S(n10936), .Z(n10077) );
  MUX2_X2 U14687 ( .A(decode_regfile_fpregs_6__9_), .B(
        decode_regfile_fpregs_7__9_), .S(n10837), .Z(n10078) );
  MUX2_X2 U14688 ( .A(decode_regfile_fpregs_4__9_), .B(
        decode_regfile_fpregs_5__9_), .S(n10837), .Z(n10079) );
  MUX2_X2 U14689 ( .A(n10079), .B(n10078), .S(n10909), .Z(n10080) );
  MUX2_X2 U14690 ( .A(decode_regfile_fpregs_2__9_), .B(
        decode_regfile_fpregs_3__9_), .S(n10837), .Z(n10081) );
  MUX2_X2 U14691 ( .A(decode_regfile_fpregs_0__9_), .B(
        decode_regfile_fpregs_1__9_), .S(n10837), .Z(n10082) );
  MUX2_X2 U14692 ( .A(n10082), .B(n10081), .S(n10909), .Z(n10083) );
  MUX2_X2 U14693 ( .A(n10083), .B(n10080), .S(n10936), .Z(n10084) );
  MUX2_X2 U14694 ( .A(n10084), .B(n10077), .S(n10950), .Z(n10085) );
  MUX2_X2 U14695 ( .A(n10085), .B(n10070), .S(n10958), .Z(decode_regfile_N50)
         );
  MUX2_X2 U14696 ( .A(decode_regfile_fpregs_30__10_), .B(
        decode_regfile_fpregs_31__10_), .S(n10838), .Z(n10086) );
  MUX2_X2 U14697 ( .A(decode_regfile_fpregs_28__10_), .B(
        decode_regfile_fpregs_29__10_), .S(n10838), .Z(n10087) );
  MUX2_X2 U14698 ( .A(n10087), .B(n10086), .S(n10910), .Z(n10088) );
  MUX2_X2 U14699 ( .A(decode_regfile_fpregs_26__10_), .B(
        decode_regfile_fpregs_27__10_), .S(n10838), .Z(n10089) );
  MUX2_X2 U14700 ( .A(decode_regfile_fpregs_24__10_), .B(
        decode_regfile_fpregs_25__10_), .S(n10838), .Z(n10090) );
  MUX2_X2 U14701 ( .A(n10090), .B(n10089), .S(n10910), .Z(n10091) );
  MUX2_X2 U14702 ( .A(n10091), .B(n10088), .S(n10937), .Z(n10092) );
  MUX2_X2 U14703 ( .A(decode_regfile_fpregs_22__10_), .B(
        decode_regfile_fpregs_23__10_), .S(n10838), .Z(n10093) );
  MUX2_X2 U14704 ( .A(decode_regfile_fpregs_20__10_), .B(
        decode_regfile_fpregs_21__10_), .S(n10838), .Z(n10094) );
  MUX2_X2 U14705 ( .A(n10094), .B(n10093), .S(n10910), .Z(n10095) );
  MUX2_X2 U14706 ( .A(decode_regfile_fpregs_18__10_), .B(
        decode_regfile_fpregs_19__10_), .S(n10838), .Z(n10096) );
  MUX2_X2 U14707 ( .A(decode_regfile_fpregs_16__10_), .B(
        decode_regfile_fpregs_17__10_), .S(n10838), .Z(n10097) );
  MUX2_X2 U14708 ( .A(n10097), .B(n10096), .S(n10910), .Z(n10098) );
  MUX2_X2 U14709 ( .A(n10098), .B(n10095), .S(n10937), .Z(n10099) );
  MUX2_X2 U14710 ( .A(n10099), .B(n10092), .S(n10951), .Z(n10100) );
  MUX2_X2 U14711 ( .A(decode_regfile_fpregs_14__10_), .B(
        decode_regfile_fpregs_15__10_), .S(n10838), .Z(n10101) );
  MUX2_X2 U14712 ( .A(decode_regfile_fpregs_12__10_), .B(
        decode_regfile_fpregs_13__10_), .S(n10838), .Z(n10102) );
  MUX2_X2 U14713 ( .A(n10102), .B(n10101), .S(n10910), .Z(n10103) );
  MUX2_X2 U14714 ( .A(decode_regfile_fpregs_10__10_), .B(
        decode_regfile_fpregs_11__10_), .S(n10838), .Z(n10104) );
  MUX2_X2 U14715 ( .A(decode_regfile_fpregs_8__10_), .B(
        decode_regfile_fpregs_9__10_), .S(n10839), .Z(n10105) );
  MUX2_X2 U14716 ( .A(n10105), .B(n10104), .S(n10910), .Z(n10106) );
  MUX2_X2 U14717 ( .A(n10106), .B(n10103), .S(n10937), .Z(n10107) );
  MUX2_X2 U14718 ( .A(decode_regfile_fpregs_6__10_), .B(
        decode_regfile_fpregs_7__10_), .S(n10839), .Z(n10108) );
  MUX2_X2 U14719 ( .A(decode_regfile_fpregs_4__10_), .B(
        decode_regfile_fpregs_5__10_), .S(n10839), .Z(n10109) );
  MUX2_X2 U14720 ( .A(n10109), .B(n10108), .S(n10910), .Z(n10110) );
  MUX2_X2 U14721 ( .A(decode_regfile_fpregs_2__10_), .B(
        decode_regfile_fpregs_3__10_), .S(n10839), .Z(n10111) );
  MUX2_X2 U14722 ( .A(decode_regfile_fpregs_0__10_), .B(
        decode_regfile_fpregs_1__10_), .S(n10839), .Z(n10112) );
  MUX2_X2 U14723 ( .A(n10112), .B(n10111), .S(n10910), .Z(n10113) );
  MUX2_X2 U14724 ( .A(n10113), .B(n10110), .S(n10937), .Z(n10114) );
  MUX2_X2 U14725 ( .A(n10114), .B(n10107), .S(n10951), .Z(n10115) );
  MUX2_X2 U14726 ( .A(n10115), .B(n10100), .S(n10959), .Z(decode_regfile_N49)
         );
  MUX2_X2 U14727 ( .A(decode_regfile_fpregs_30__11_), .B(
        decode_regfile_fpregs_31__11_), .S(n10839), .Z(n10116) );
  MUX2_X2 U14728 ( .A(decode_regfile_fpregs_28__11_), .B(
        decode_regfile_fpregs_29__11_), .S(n10839), .Z(n10117) );
  MUX2_X2 U14729 ( .A(n10117), .B(n10116), .S(n10910), .Z(n10118) );
  MUX2_X2 U14730 ( .A(decode_regfile_fpregs_26__11_), .B(
        decode_regfile_fpregs_27__11_), .S(n10839), .Z(n10119) );
  MUX2_X2 U14731 ( .A(decode_regfile_fpregs_24__11_), .B(
        decode_regfile_fpregs_25__11_), .S(n10839), .Z(n10120) );
  MUX2_X2 U14732 ( .A(n10120), .B(n10119), .S(n10910), .Z(n10121) );
  MUX2_X2 U14733 ( .A(n10121), .B(n10118), .S(n10937), .Z(n10122) );
  MUX2_X2 U14734 ( .A(decode_regfile_fpregs_22__11_), .B(
        decode_regfile_fpregs_23__11_), .S(n10839), .Z(n10123) );
  MUX2_X2 U14735 ( .A(decode_regfile_fpregs_20__11_), .B(
        decode_regfile_fpregs_21__11_), .S(n10839), .Z(n10124) );
  MUX2_X2 U14736 ( .A(n10124), .B(n10123), .S(n10910), .Z(n10125) );
  MUX2_X2 U14737 ( .A(decode_regfile_fpregs_18__11_), .B(
        decode_regfile_fpregs_19__11_), .S(n10840), .Z(n10126) );
  MUX2_X2 U14738 ( .A(decode_regfile_fpregs_16__11_), .B(
        decode_regfile_fpregs_17__11_), .S(n10840), .Z(n10127) );
  MUX2_X2 U14739 ( .A(n10127), .B(n10126), .S(n10911), .Z(n10128) );
  MUX2_X2 U14740 ( .A(n10128), .B(n10125), .S(n10937), .Z(n10129) );
  MUX2_X2 U14741 ( .A(n10129), .B(n10122), .S(n10951), .Z(n10130) );
  MUX2_X2 U14742 ( .A(decode_regfile_fpregs_14__11_), .B(
        decode_regfile_fpregs_15__11_), .S(n10840), .Z(n10131) );
  MUX2_X2 U14743 ( .A(decode_regfile_fpregs_12__11_), .B(
        decode_regfile_fpregs_13__11_), .S(n10840), .Z(n10132) );
  MUX2_X2 U14744 ( .A(n10132), .B(n10131), .S(n10911), .Z(n10133) );
  MUX2_X2 U14745 ( .A(decode_regfile_fpregs_10__11_), .B(
        decode_regfile_fpregs_11__11_), .S(n10840), .Z(n10134) );
  MUX2_X2 U14746 ( .A(decode_regfile_fpregs_8__11_), .B(
        decode_regfile_fpregs_9__11_), .S(n10840), .Z(n10135) );
  MUX2_X2 U14747 ( .A(n10135), .B(n10134), .S(n10911), .Z(n10136) );
  MUX2_X2 U14748 ( .A(n10136), .B(n10133), .S(n10937), .Z(n10137) );
  MUX2_X2 U14749 ( .A(decode_regfile_fpregs_6__11_), .B(
        decode_regfile_fpregs_7__11_), .S(n10840), .Z(n10138) );
  MUX2_X2 U14750 ( .A(decode_regfile_fpregs_4__11_), .B(
        decode_regfile_fpregs_5__11_), .S(n10840), .Z(n10139) );
  MUX2_X2 U14751 ( .A(n10139), .B(n10138), .S(n10911), .Z(n10140) );
  MUX2_X2 U14752 ( .A(decode_regfile_fpregs_2__11_), .B(
        decode_regfile_fpregs_3__11_), .S(n10840), .Z(n10141) );
  MUX2_X2 U14753 ( .A(decode_regfile_fpregs_0__11_), .B(
        decode_regfile_fpregs_1__11_), .S(n10840), .Z(n10142) );
  MUX2_X2 U14754 ( .A(n10142), .B(n10141), .S(n10911), .Z(n10143) );
  MUX2_X2 U14755 ( .A(n10143), .B(n10140), .S(n10937), .Z(n10144) );
  MUX2_X2 U14756 ( .A(n10144), .B(n10137), .S(n10951), .Z(n10145) );
  MUX2_X2 U14757 ( .A(n10145), .B(n10130), .S(n10959), .Z(decode_regfile_N48)
         );
  MUX2_X2 U14758 ( .A(decode_regfile_fpregs_30__12_), .B(
        decode_regfile_fpregs_31__12_), .S(n10840), .Z(n10146) );
  MUX2_X2 U14759 ( .A(decode_regfile_fpregs_28__12_), .B(
        decode_regfile_fpregs_29__12_), .S(n10841), .Z(n10147) );
  MUX2_X2 U14760 ( .A(n10147), .B(n10146), .S(n10911), .Z(n10148) );
  MUX2_X2 U14761 ( .A(decode_regfile_fpregs_26__12_), .B(
        decode_regfile_fpregs_27__12_), .S(n10841), .Z(n10149) );
  MUX2_X2 U14762 ( .A(decode_regfile_fpregs_24__12_), .B(
        decode_regfile_fpregs_25__12_), .S(n10841), .Z(n10150) );
  MUX2_X2 U14763 ( .A(n10150), .B(n10149), .S(n10911), .Z(n10151) );
  MUX2_X2 U14764 ( .A(n10151), .B(n10148), .S(n10937), .Z(n10152) );
  MUX2_X2 U14765 ( .A(decode_regfile_fpregs_22__12_), .B(
        decode_regfile_fpregs_23__12_), .S(n10841), .Z(n10153) );
  MUX2_X2 U14766 ( .A(decode_regfile_fpregs_20__12_), .B(
        decode_regfile_fpregs_21__12_), .S(n10841), .Z(n10154) );
  MUX2_X2 U14767 ( .A(n10154), .B(n10153), .S(n10911), .Z(n10155) );
  MUX2_X2 U14768 ( .A(decode_regfile_fpregs_18__12_), .B(
        decode_regfile_fpregs_19__12_), .S(n10841), .Z(n10156) );
  MUX2_X2 U14769 ( .A(decode_regfile_fpregs_16__12_), .B(
        decode_regfile_fpregs_17__12_), .S(n10841), .Z(n10157) );
  MUX2_X2 U14770 ( .A(n10157), .B(n10156), .S(n10911), .Z(n10158) );
  MUX2_X2 U14771 ( .A(n10158), .B(n10155), .S(n10937), .Z(n10159) );
  MUX2_X2 U14772 ( .A(n10159), .B(n10152), .S(n10951), .Z(n10160) );
  MUX2_X2 U14773 ( .A(decode_regfile_fpregs_14__12_), .B(
        decode_regfile_fpregs_15__12_), .S(n10841), .Z(n10161) );
  MUX2_X2 U14774 ( .A(decode_regfile_fpregs_12__12_), .B(
        decode_regfile_fpregs_13__12_), .S(n10841), .Z(n10162) );
  MUX2_X2 U14775 ( .A(n10162), .B(n10161), .S(n10911), .Z(n10163) );
  MUX2_X2 U14776 ( .A(decode_regfile_fpregs_10__12_), .B(
        decode_regfile_fpregs_11__12_), .S(n10841), .Z(n10164) );
  MUX2_X2 U14777 ( .A(decode_regfile_fpregs_8__12_), .B(
        decode_regfile_fpregs_9__12_), .S(n10841), .Z(n10165) );
  MUX2_X2 U14778 ( .A(n10165), .B(n10164), .S(n10911), .Z(n10166) );
  MUX2_X2 U14779 ( .A(n10166), .B(n10163), .S(n10937), .Z(n10167) );
  MUX2_X2 U14780 ( .A(decode_regfile_fpregs_6__12_), .B(
        decode_regfile_fpregs_7__12_), .S(n10842), .Z(n10168) );
  MUX2_X2 U14781 ( .A(decode_regfile_fpregs_4__12_), .B(
        decode_regfile_fpregs_5__12_), .S(n10842), .Z(n10169) );
  MUX2_X2 U14782 ( .A(n10169), .B(n10168), .S(n10912), .Z(n10170) );
  MUX2_X2 U14783 ( .A(decode_regfile_fpregs_2__12_), .B(
        decode_regfile_fpregs_3__12_), .S(n10842), .Z(n10171) );
  MUX2_X2 U14784 ( .A(decode_regfile_fpregs_0__12_), .B(
        decode_regfile_fpregs_1__12_), .S(n10842), .Z(n10172) );
  MUX2_X2 U14785 ( .A(n10172), .B(n10171), .S(n10912), .Z(n10173) );
  MUX2_X2 U14786 ( .A(n10173), .B(n10170), .S(n10938), .Z(n10174) );
  MUX2_X2 U14787 ( .A(n10174), .B(n10167), .S(n10951), .Z(n10175) );
  MUX2_X2 U14788 ( .A(n10175), .B(n10160), .S(n10959), .Z(decode_regfile_N47)
         );
  MUX2_X2 U14789 ( .A(decode_regfile_fpregs_30__13_), .B(
        decode_regfile_fpregs_31__13_), .S(n10842), .Z(n10176) );
  MUX2_X2 U14790 ( .A(decode_regfile_fpregs_28__13_), .B(
        decode_regfile_fpregs_29__13_), .S(n10842), .Z(n10177) );
  MUX2_X2 U14791 ( .A(n10177), .B(n10176), .S(n10912), .Z(n10178) );
  MUX2_X2 U14792 ( .A(decode_regfile_fpregs_26__13_), .B(
        decode_regfile_fpregs_27__13_), .S(n10842), .Z(n10179) );
  MUX2_X2 U14793 ( .A(decode_regfile_fpregs_24__13_), .B(
        decode_regfile_fpregs_25__13_), .S(n10842), .Z(n10180) );
  MUX2_X2 U14794 ( .A(n10180), .B(n10179), .S(n10912), .Z(n10181) );
  MUX2_X2 U14795 ( .A(n10181), .B(n10178), .S(n10938), .Z(n10182) );
  MUX2_X2 U14796 ( .A(decode_regfile_fpregs_22__13_), .B(
        decode_regfile_fpregs_23__13_), .S(n10842), .Z(n10183) );
  MUX2_X2 U14797 ( .A(decode_regfile_fpregs_20__13_), .B(
        decode_regfile_fpregs_21__13_), .S(n10842), .Z(n10184) );
  MUX2_X2 U14798 ( .A(n10184), .B(n10183), .S(n10912), .Z(n10185) );
  MUX2_X2 U14799 ( .A(decode_regfile_fpregs_18__13_), .B(
        decode_regfile_fpregs_19__13_), .S(n10842), .Z(n10186) );
  MUX2_X2 U14800 ( .A(decode_regfile_fpregs_16__13_), .B(
        decode_regfile_fpregs_17__13_), .S(n10843), .Z(n10187) );
  MUX2_X2 U14801 ( .A(n10187), .B(n10186), .S(n10912), .Z(n10188) );
  MUX2_X2 U14802 ( .A(n10188), .B(n10185), .S(n10938), .Z(n10189) );
  MUX2_X2 U14803 ( .A(n10189), .B(n10182), .S(n10951), .Z(n10190) );
  MUX2_X2 U14804 ( .A(decode_regfile_fpregs_14__13_), .B(
        decode_regfile_fpregs_15__13_), .S(n10843), .Z(n10191) );
  MUX2_X2 U14805 ( .A(decode_regfile_fpregs_12__13_), .B(
        decode_regfile_fpregs_13__13_), .S(n10843), .Z(n10192) );
  MUX2_X2 U14806 ( .A(n10192), .B(n10191), .S(n10912), .Z(n10193) );
  MUX2_X2 U14807 ( .A(decode_regfile_fpregs_10__13_), .B(
        decode_regfile_fpregs_11__13_), .S(n10843), .Z(n10194) );
  MUX2_X2 U14808 ( .A(decode_regfile_fpregs_8__13_), .B(
        decode_regfile_fpregs_9__13_), .S(n10843), .Z(n10195) );
  MUX2_X2 U14809 ( .A(n10195), .B(n10194), .S(n10912), .Z(n10196) );
  MUX2_X2 U14810 ( .A(n10196), .B(n10193), .S(n10938), .Z(n10197) );
  MUX2_X2 U14811 ( .A(decode_regfile_fpregs_6__13_), .B(
        decode_regfile_fpregs_7__13_), .S(n10843), .Z(n10198) );
  MUX2_X2 U14812 ( .A(decode_regfile_fpregs_4__13_), .B(
        decode_regfile_fpregs_5__13_), .S(n10843), .Z(n10199) );
  MUX2_X2 U14813 ( .A(n10199), .B(n10198), .S(n10912), .Z(n10200) );
  MUX2_X2 U14814 ( .A(decode_regfile_fpregs_2__13_), .B(
        decode_regfile_fpregs_3__13_), .S(n10843), .Z(n10201) );
  MUX2_X2 U14815 ( .A(decode_regfile_fpregs_0__13_), .B(
        decode_regfile_fpregs_1__13_), .S(n10843), .Z(n10202) );
  MUX2_X2 U14816 ( .A(n10202), .B(n10201), .S(n10912), .Z(n10203) );
  MUX2_X2 U14817 ( .A(n10203), .B(n10200), .S(n10938), .Z(n10204) );
  MUX2_X2 U14818 ( .A(n10204), .B(n10197), .S(n10951), .Z(n10205) );
  MUX2_X2 U14819 ( .A(n10205), .B(n10190), .S(n10959), .Z(decode_regfile_N46)
         );
  MUX2_X2 U14820 ( .A(decode_regfile_fpregs_30__14_), .B(
        decode_regfile_fpregs_31__14_), .S(n10843), .Z(n10206) );
  MUX2_X2 U14821 ( .A(decode_regfile_fpregs_28__14_), .B(
        decode_regfile_fpregs_29__14_), .S(n10843), .Z(n10207) );
  MUX2_X2 U14822 ( .A(n10207), .B(n10206), .S(n10912), .Z(n10208) );
  MUX2_X2 U14823 ( .A(decode_regfile_fpregs_26__14_), .B(
        decode_regfile_fpregs_27__14_), .S(n10844), .Z(n10209) );
  MUX2_X2 U14824 ( .A(decode_regfile_fpregs_24__14_), .B(
        decode_regfile_fpregs_25__14_), .S(n10844), .Z(n10210) );
  MUX2_X2 U14825 ( .A(n10210), .B(n10209), .S(n10913), .Z(n10211) );
  MUX2_X2 U14826 ( .A(n10211), .B(n10208), .S(n10938), .Z(n10212) );
  MUX2_X2 U14827 ( .A(decode_regfile_fpregs_22__14_), .B(
        decode_regfile_fpregs_23__14_), .S(n10844), .Z(n10213) );
  MUX2_X2 U14828 ( .A(decode_regfile_fpregs_20__14_), .B(
        decode_regfile_fpregs_21__14_), .S(n10844), .Z(n10214) );
  MUX2_X2 U14829 ( .A(n10214), .B(n10213), .S(n10913), .Z(n10215) );
  MUX2_X2 U14830 ( .A(decode_regfile_fpregs_18__14_), .B(
        decode_regfile_fpregs_19__14_), .S(n10844), .Z(n10216) );
  MUX2_X2 U14831 ( .A(decode_regfile_fpregs_16__14_), .B(
        decode_regfile_fpregs_17__14_), .S(n10844), .Z(n10217) );
  MUX2_X2 U14832 ( .A(n10217), .B(n10216), .S(n10913), .Z(n10218) );
  MUX2_X2 U14833 ( .A(n10218), .B(n10215), .S(n10938), .Z(n10219) );
  MUX2_X2 U14834 ( .A(n10219), .B(n10212), .S(n10951), .Z(n10220) );
  MUX2_X2 U14835 ( .A(decode_regfile_fpregs_14__14_), .B(
        decode_regfile_fpregs_15__14_), .S(n10844), .Z(n10221) );
  MUX2_X2 U14836 ( .A(decode_regfile_fpregs_12__14_), .B(
        decode_regfile_fpregs_13__14_), .S(n10844), .Z(n10222) );
  MUX2_X2 U14837 ( .A(n10222), .B(n10221), .S(n10913), .Z(n10223) );
  MUX2_X2 U14838 ( .A(decode_regfile_fpregs_10__14_), .B(
        decode_regfile_fpregs_11__14_), .S(n10844), .Z(n10224) );
  MUX2_X2 U14839 ( .A(decode_regfile_fpregs_8__14_), .B(
        decode_regfile_fpregs_9__14_), .S(n10844), .Z(n10225) );
  MUX2_X2 U14840 ( .A(n10225), .B(n10224), .S(n10913), .Z(n10226) );
  MUX2_X2 U14841 ( .A(n10226), .B(n10223), .S(n10938), .Z(n10227) );
  MUX2_X2 U14842 ( .A(decode_regfile_fpregs_6__14_), .B(
        decode_regfile_fpregs_7__14_), .S(n10844), .Z(n10228) );
  MUX2_X2 U14843 ( .A(decode_regfile_fpregs_4__14_), .B(
        decode_regfile_fpregs_5__14_), .S(n10845), .Z(n10229) );
  MUX2_X2 U14844 ( .A(n10229), .B(n10228), .S(n10913), .Z(n10230) );
  MUX2_X2 U14845 ( .A(decode_regfile_fpregs_2__14_), .B(
        decode_regfile_fpregs_3__14_), .S(n10845), .Z(n10231) );
  MUX2_X2 U14846 ( .A(decode_regfile_fpregs_0__14_), .B(
        decode_regfile_fpregs_1__14_), .S(n10845), .Z(n10232) );
  MUX2_X2 U14847 ( .A(n10232), .B(n10231), .S(n10913), .Z(n10233) );
  MUX2_X2 U14848 ( .A(n10233), .B(n10230), .S(n10938), .Z(n10234) );
  MUX2_X2 U14849 ( .A(n10234), .B(n10227), .S(n10951), .Z(n10235) );
  MUX2_X2 U14850 ( .A(n10235), .B(n10220), .S(n10959), .Z(decode_regfile_N45)
         );
  MUX2_X2 U14851 ( .A(decode_regfile_fpregs_30__15_), .B(
        decode_regfile_fpregs_31__15_), .S(n10845), .Z(n10236) );
  MUX2_X2 U14852 ( .A(decode_regfile_fpregs_28__15_), .B(
        decode_regfile_fpregs_29__15_), .S(n10845), .Z(n10237) );
  MUX2_X2 U14853 ( .A(n10237), .B(n10236), .S(n10913), .Z(n10238) );
  MUX2_X2 U14854 ( .A(decode_regfile_fpregs_26__15_), .B(
        decode_regfile_fpregs_27__15_), .S(n10845), .Z(n10239) );
  MUX2_X2 U14855 ( .A(decode_regfile_fpregs_24__15_), .B(
        decode_regfile_fpregs_25__15_), .S(n10845), .Z(n10240) );
  MUX2_X2 U14856 ( .A(n10240), .B(n10239), .S(n10913), .Z(n10241) );
  MUX2_X2 U14857 ( .A(n10241), .B(n10238), .S(n10938), .Z(n10242) );
  MUX2_X2 U14858 ( .A(decode_regfile_fpregs_22__15_), .B(
        decode_regfile_fpregs_23__15_), .S(n10845), .Z(n10243) );
  MUX2_X2 U14859 ( .A(decode_regfile_fpregs_20__15_), .B(
        decode_regfile_fpregs_21__15_), .S(n10845), .Z(n10244) );
  MUX2_X2 U14860 ( .A(n10244), .B(n10243), .S(n10913), .Z(n10245) );
  MUX2_X2 U14861 ( .A(decode_regfile_fpregs_18__15_), .B(
        decode_regfile_fpregs_19__15_), .S(n10845), .Z(n10246) );
  MUX2_X2 U14862 ( .A(decode_regfile_fpregs_16__15_), .B(
        decode_regfile_fpregs_17__15_), .S(n10845), .Z(n10247) );
  MUX2_X2 U14863 ( .A(n10247), .B(n10246), .S(n10913), .Z(n10248) );
  MUX2_X2 U14864 ( .A(n10248), .B(n10245), .S(n10938), .Z(n10249) );
  MUX2_X2 U14865 ( .A(n10249), .B(n10242), .S(n10951), .Z(n10250) );
  MUX2_X2 U14866 ( .A(decode_regfile_fpregs_14__15_), .B(
        decode_regfile_fpregs_15__15_), .S(n10846), .Z(n10251) );
  MUX2_X2 U14867 ( .A(decode_regfile_fpregs_12__15_), .B(
        decode_regfile_fpregs_13__15_), .S(n10846), .Z(n10252) );
  MUX2_X2 U14868 ( .A(n10252), .B(n10251), .S(n10914), .Z(n10253) );
  MUX2_X2 U14869 ( .A(decode_regfile_fpregs_10__15_), .B(
        decode_regfile_fpregs_11__15_), .S(n10846), .Z(n10254) );
  MUX2_X2 U14870 ( .A(decode_regfile_fpregs_8__15_), .B(
        decode_regfile_fpregs_9__15_), .S(n10846), .Z(n10255) );
  MUX2_X2 U14871 ( .A(n10255), .B(n10254), .S(n10914), .Z(n10256) );
  MUX2_X2 U14872 ( .A(n10256), .B(n10253), .S(n10939), .Z(n10257) );
  MUX2_X2 U14873 ( .A(decode_regfile_fpregs_6__15_), .B(
        decode_regfile_fpregs_7__15_), .S(n10846), .Z(n10258) );
  MUX2_X2 U14874 ( .A(decode_regfile_fpregs_4__15_), .B(
        decode_regfile_fpregs_5__15_), .S(n10846), .Z(n10259) );
  MUX2_X2 U14875 ( .A(n10259), .B(n10258), .S(n10914), .Z(n10260) );
  MUX2_X2 U14876 ( .A(decode_regfile_fpregs_2__15_), .B(
        decode_regfile_fpregs_3__15_), .S(n10846), .Z(n10261) );
  MUX2_X2 U14877 ( .A(decode_regfile_fpregs_0__15_), .B(
        decode_regfile_fpregs_1__15_), .S(n10846), .Z(n10262) );
  MUX2_X2 U14878 ( .A(n10262), .B(n10261), .S(n10914), .Z(n10263) );
  MUX2_X2 U14879 ( .A(n10263), .B(n10260), .S(n10939), .Z(n10264) );
  MUX2_X2 U14880 ( .A(n10264), .B(n10257), .S(n10952), .Z(n10265) );
  MUX2_X2 U14881 ( .A(n10265), .B(n10250), .S(n10959), .Z(decode_regfile_N44)
         );
  MUX2_X2 U14882 ( .A(decode_regfile_fpregs_30__16_), .B(
        decode_regfile_fpregs_31__16_), .S(n10846), .Z(n10266) );
  MUX2_X2 U14883 ( .A(decode_regfile_fpregs_28__16_), .B(
        decode_regfile_fpregs_29__16_), .S(n10846), .Z(n10267) );
  MUX2_X2 U14884 ( .A(n10267), .B(n10266), .S(n10914), .Z(n10268) );
  MUX2_X2 U14885 ( .A(decode_regfile_fpregs_26__16_), .B(
        decode_regfile_fpregs_27__16_), .S(n10846), .Z(n10269) );
  MUX2_X2 U14886 ( .A(decode_regfile_fpregs_24__16_), .B(
        decode_regfile_fpregs_25__16_), .S(n10847), .Z(n10270) );
  MUX2_X2 U14887 ( .A(n10270), .B(n10269), .S(n10914), .Z(n10271) );
  MUX2_X2 U14888 ( .A(n10271), .B(n10268), .S(n10939), .Z(n10272) );
  MUX2_X2 U14889 ( .A(decode_regfile_fpregs_22__16_), .B(
        decode_regfile_fpregs_23__16_), .S(n10847), .Z(n10273) );
  MUX2_X2 U14890 ( .A(decode_regfile_fpregs_20__16_), .B(
        decode_regfile_fpregs_21__16_), .S(n10847), .Z(n10274) );
  MUX2_X2 U14891 ( .A(n10274), .B(n10273), .S(n10914), .Z(n10275) );
  MUX2_X2 U14892 ( .A(decode_regfile_fpregs_18__16_), .B(
        decode_regfile_fpregs_19__16_), .S(n10847), .Z(n10276) );
  MUX2_X2 U14893 ( .A(decode_regfile_fpregs_16__16_), .B(
        decode_regfile_fpregs_17__16_), .S(n10847), .Z(n10277) );
  MUX2_X2 U14894 ( .A(n10277), .B(n10276), .S(n10914), .Z(n10278) );
  MUX2_X2 U14895 ( .A(n10278), .B(n10275), .S(n10939), .Z(n10279) );
  MUX2_X2 U14896 ( .A(n10279), .B(n10272), .S(n10952), .Z(n10280) );
  MUX2_X2 U14897 ( .A(decode_regfile_fpregs_14__16_), .B(
        decode_regfile_fpregs_15__16_), .S(n10847), .Z(n10281) );
  MUX2_X2 U14898 ( .A(decode_regfile_fpregs_12__16_), .B(
        decode_regfile_fpregs_13__16_), .S(n10847), .Z(n10282) );
  MUX2_X2 U14899 ( .A(n10282), .B(n10281), .S(n10914), .Z(n10283) );
  MUX2_X2 U14900 ( .A(decode_regfile_fpregs_10__16_), .B(
        decode_regfile_fpregs_11__16_), .S(n10847), .Z(n10284) );
  MUX2_X2 U14901 ( .A(decode_regfile_fpregs_8__16_), .B(
        decode_regfile_fpregs_9__16_), .S(n10847), .Z(n10285) );
  MUX2_X2 U14902 ( .A(n10285), .B(n10284), .S(n10914), .Z(n10286) );
  MUX2_X2 U14903 ( .A(n10286), .B(n10283), .S(n10939), .Z(n10287) );
  MUX2_X2 U14904 ( .A(decode_regfile_fpregs_6__16_), .B(
        decode_regfile_fpregs_7__16_), .S(n10847), .Z(n10288) );
  MUX2_X2 U14905 ( .A(decode_regfile_fpregs_4__16_), .B(
        decode_regfile_fpregs_5__16_), .S(n10847), .Z(n10289) );
  MUX2_X2 U14906 ( .A(n10289), .B(n10288), .S(n10914), .Z(n10290) );
  MUX2_X2 U14907 ( .A(decode_regfile_fpregs_2__16_), .B(
        decode_regfile_fpregs_3__16_), .S(n10848), .Z(n10291) );
  MUX2_X2 U14908 ( .A(decode_regfile_fpregs_0__16_), .B(
        decode_regfile_fpregs_1__16_), .S(n10848), .Z(n10292) );
  MUX2_X2 U14909 ( .A(n10292), .B(n10291), .S(n10915), .Z(n10293) );
  MUX2_X2 U14910 ( .A(n10293), .B(n10290), .S(n10939), .Z(n10294) );
  MUX2_X2 U14911 ( .A(n10294), .B(n10287), .S(n10952), .Z(n10295) );
  MUX2_X2 U14912 ( .A(n10295), .B(n10280), .S(n10959), .Z(decode_regfile_N43)
         );
  MUX2_X2 U14913 ( .A(decode_regfile_fpregs_30__17_), .B(
        decode_regfile_fpregs_31__17_), .S(n10848), .Z(n10296) );
  MUX2_X2 U14914 ( .A(decode_regfile_fpregs_28__17_), .B(
        decode_regfile_fpregs_29__17_), .S(n10848), .Z(n10297) );
  MUX2_X2 U14915 ( .A(n10297), .B(n10296), .S(n10915), .Z(n10298) );
  MUX2_X2 U14916 ( .A(decode_regfile_fpregs_26__17_), .B(
        decode_regfile_fpregs_27__17_), .S(n10848), .Z(n10299) );
  MUX2_X2 U14917 ( .A(decode_regfile_fpregs_24__17_), .B(
        decode_regfile_fpregs_25__17_), .S(n10848), .Z(n10300) );
  MUX2_X2 U14918 ( .A(n10300), .B(n10299), .S(n10915), .Z(n10301) );
  MUX2_X2 U14919 ( .A(n10301), .B(n10298), .S(n10939), .Z(n10302) );
  MUX2_X2 U14920 ( .A(decode_regfile_fpregs_22__17_), .B(
        decode_regfile_fpregs_23__17_), .S(n10848), .Z(n10303) );
  MUX2_X2 U14921 ( .A(decode_regfile_fpregs_20__17_), .B(
        decode_regfile_fpregs_21__17_), .S(n10848), .Z(n10304) );
  MUX2_X2 U14922 ( .A(n10304), .B(n10303), .S(n10915), .Z(n10305) );
  MUX2_X2 U14923 ( .A(decode_regfile_fpregs_18__17_), .B(
        decode_regfile_fpregs_19__17_), .S(n10848), .Z(n10306) );
  MUX2_X2 U14924 ( .A(decode_regfile_fpregs_16__17_), .B(
        decode_regfile_fpregs_17__17_), .S(n10848), .Z(n10307) );
  MUX2_X2 U14925 ( .A(n10307), .B(n10306), .S(n10915), .Z(n10308) );
  MUX2_X2 U14926 ( .A(n10308), .B(n10305), .S(n10939), .Z(n10309) );
  MUX2_X2 U14927 ( .A(n10309), .B(n10302), .S(n10952), .Z(n10310) );
  MUX2_X2 U14928 ( .A(decode_regfile_fpregs_14__17_), .B(
        decode_regfile_fpregs_15__17_), .S(n10848), .Z(n10311) );
  MUX2_X2 U14929 ( .A(decode_regfile_fpregs_12__17_), .B(
        decode_regfile_fpregs_13__17_), .S(n10849), .Z(n10312) );
  MUX2_X2 U14930 ( .A(n10312), .B(n10311), .S(n10915), .Z(n10313) );
  MUX2_X2 U14931 ( .A(decode_regfile_fpregs_10__17_), .B(
        decode_regfile_fpregs_11__17_), .S(n10849), .Z(n10314) );
  MUX2_X2 U14932 ( .A(decode_regfile_fpregs_8__17_), .B(
        decode_regfile_fpregs_9__17_), .S(n10849), .Z(n10315) );
  MUX2_X2 U14933 ( .A(n10315), .B(n10314), .S(n10915), .Z(n10316) );
  MUX2_X2 U14934 ( .A(n10316), .B(n10313), .S(n10939), .Z(n10317) );
  MUX2_X2 U14935 ( .A(decode_regfile_fpregs_6__17_), .B(
        decode_regfile_fpregs_7__17_), .S(n10849), .Z(n10318) );
  MUX2_X2 U14936 ( .A(decode_regfile_fpregs_4__17_), .B(
        decode_regfile_fpregs_5__17_), .S(n10849), .Z(n10319) );
  MUX2_X2 U14937 ( .A(n10319), .B(n10318), .S(n10915), .Z(n10320) );
  MUX2_X2 U14938 ( .A(decode_regfile_fpregs_2__17_), .B(
        decode_regfile_fpregs_3__17_), .S(n10849), .Z(n10321) );
  MUX2_X2 U14939 ( .A(decode_regfile_fpregs_0__17_), .B(
        decode_regfile_fpregs_1__17_), .S(n10849), .Z(n10322) );
  MUX2_X2 U14940 ( .A(n10322), .B(n10321), .S(n10915), .Z(n10323) );
  MUX2_X2 U14941 ( .A(n10323), .B(n10320), .S(n10939), .Z(n10324) );
  MUX2_X2 U14942 ( .A(n10324), .B(n10317), .S(n10952), .Z(n10325) );
  MUX2_X2 U14943 ( .A(n10325), .B(n10310), .S(n10959), .Z(decode_regfile_N42)
         );
  MUX2_X2 U14944 ( .A(decode_regfile_fpregs_30__18_), .B(
        decode_regfile_fpregs_31__18_), .S(n10849), .Z(n10326) );
  MUX2_X2 U14945 ( .A(decode_regfile_fpregs_28__18_), .B(
        decode_regfile_fpregs_29__18_), .S(n10849), .Z(n10327) );
  MUX2_X2 U14946 ( .A(n10327), .B(n10326), .S(n10915), .Z(n10328) );
  MUX2_X2 U14947 ( .A(decode_regfile_fpregs_26__18_), .B(
        decode_regfile_fpregs_27__18_), .S(n10849), .Z(n10329) );
  MUX2_X2 U14948 ( .A(decode_regfile_fpregs_24__18_), .B(
        decode_regfile_fpregs_25__18_), .S(n10849), .Z(n10330) );
  MUX2_X2 U14949 ( .A(n10330), .B(n10329), .S(n10915), .Z(n10331) );
  MUX2_X2 U14950 ( .A(n10331), .B(n10328), .S(n10939), .Z(n10332) );
  MUX2_X2 U14951 ( .A(decode_regfile_fpregs_22__18_), .B(
        decode_regfile_fpregs_23__18_), .S(n10850), .Z(n10333) );
  MUX2_X2 U14952 ( .A(decode_regfile_fpregs_20__18_), .B(
        decode_regfile_fpregs_21__18_), .S(n10850), .Z(n10334) );
  MUX2_X2 U14953 ( .A(n10334), .B(n10333), .S(n10916), .Z(n10335) );
  MUX2_X2 U14954 ( .A(decode_regfile_fpregs_18__18_), .B(
        decode_regfile_fpregs_19__18_), .S(n10850), .Z(n10336) );
  MUX2_X2 U14955 ( .A(decode_regfile_fpregs_16__18_), .B(
        decode_regfile_fpregs_17__18_), .S(n10850), .Z(n10337) );
  MUX2_X2 U14956 ( .A(n10337), .B(n10336), .S(n10916), .Z(n10338) );
  MUX2_X2 U14957 ( .A(n10338), .B(n10335), .S(n10940), .Z(n10339) );
  MUX2_X2 U14958 ( .A(n10339), .B(n10332), .S(n10952), .Z(n10340) );
  MUX2_X2 U14959 ( .A(decode_regfile_fpregs_14__18_), .B(
        decode_regfile_fpregs_15__18_), .S(n10850), .Z(n10341) );
  MUX2_X2 U14960 ( .A(decode_regfile_fpregs_12__18_), .B(
        decode_regfile_fpregs_13__18_), .S(n10850), .Z(n10342) );
  MUX2_X2 U14961 ( .A(n10342), .B(n10341), .S(n10916), .Z(n10343) );
  MUX2_X2 U14962 ( .A(decode_regfile_fpregs_10__18_), .B(
        decode_regfile_fpregs_11__18_), .S(n10850), .Z(n10344) );
  MUX2_X2 U14963 ( .A(decode_regfile_fpregs_8__18_), .B(
        decode_regfile_fpregs_9__18_), .S(n10850), .Z(n10345) );
  MUX2_X2 U14964 ( .A(n10345), .B(n10344), .S(n10916), .Z(n10346) );
  MUX2_X2 U14965 ( .A(n10346), .B(n10343), .S(n10940), .Z(n10347) );
  MUX2_X2 U14966 ( .A(decode_regfile_fpregs_6__18_), .B(
        decode_regfile_fpregs_7__18_), .S(n10850), .Z(n10348) );
  MUX2_X2 U14967 ( .A(decode_regfile_fpregs_4__18_), .B(
        decode_regfile_fpregs_5__18_), .S(n10850), .Z(n10349) );
  MUX2_X2 U14968 ( .A(n10349), .B(n10348), .S(n10916), .Z(n10350) );
  MUX2_X2 U14969 ( .A(decode_regfile_fpregs_2__18_), .B(
        decode_regfile_fpregs_3__18_), .S(n10850), .Z(n10351) );
  MUX2_X2 U14970 ( .A(decode_regfile_fpregs_0__18_), .B(
        decode_regfile_fpregs_1__18_), .S(n10851), .Z(n10352) );
  MUX2_X2 U14971 ( .A(n10352), .B(n10351), .S(n10916), .Z(n10353) );
  MUX2_X2 U14972 ( .A(n10353), .B(n10350), .S(n10940), .Z(n10354) );
  MUX2_X2 U14973 ( .A(n10354), .B(n10347), .S(n10952), .Z(n10355) );
  MUX2_X2 U14974 ( .A(n10355), .B(n10340), .S(n10959), .Z(decode_regfile_N41)
         );
  MUX2_X2 U14975 ( .A(decode_regfile_fpregs_30__19_), .B(
        decode_regfile_fpregs_31__19_), .S(n10851), .Z(n10356) );
  MUX2_X2 U14976 ( .A(decode_regfile_fpregs_28__19_), .B(
        decode_regfile_fpregs_29__19_), .S(n10851), .Z(n10357) );
  MUX2_X2 U14977 ( .A(n10357), .B(n10356), .S(n10916), .Z(n10358) );
  MUX2_X2 U14978 ( .A(decode_regfile_fpregs_26__19_), .B(
        decode_regfile_fpregs_27__19_), .S(n10851), .Z(n10359) );
  MUX2_X2 U14979 ( .A(decode_regfile_fpregs_24__19_), .B(
        decode_regfile_fpregs_25__19_), .S(n10851), .Z(n10360) );
  MUX2_X2 U14980 ( .A(n10360), .B(n10359), .S(n10916), .Z(n10361) );
  MUX2_X2 U14981 ( .A(n10361), .B(n10358), .S(n10940), .Z(n10362) );
  MUX2_X2 U14982 ( .A(decode_regfile_fpregs_22__19_), .B(
        decode_regfile_fpregs_23__19_), .S(n10851), .Z(n10363) );
  MUX2_X2 U14983 ( .A(decode_regfile_fpregs_20__19_), .B(
        decode_regfile_fpregs_21__19_), .S(n10851), .Z(n10364) );
  MUX2_X2 U14984 ( .A(n10364), .B(n10363), .S(n10916), .Z(n10365) );
  MUX2_X2 U14985 ( .A(decode_regfile_fpregs_18__19_), .B(
        decode_regfile_fpregs_19__19_), .S(n10851), .Z(n10366) );
  MUX2_X2 U14986 ( .A(decode_regfile_fpregs_16__19_), .B(
        decode_regfile_fpregs_17__19_), .S(n10851), .Z(n10367) );
  MUX2_X2 U14987 ( .A(n10367), .B(n10366), .S(n10916), .Z(n10368) );
  MUX2_X2 U14988 ( .A(n10368), .B(n10365), .S(n10940), .Z(n10369) );
  MUX2_X2 U14989 ( .A(n10369), .B(n10362), .S(n10952), .Z(n10370) );
  MUX2_X2 U14990 ( .A(decode_regfile_fpregs_14__19_), .B(
        decode_regfile_fpregs_15__19_), .S(n10851), .Z(n10371) );
  MUX2_X2 U14991 ( .A(decode_regfile_fpregs_12__19_), .B(
        decode_regfile_fpregs_13__19_), .S(n10851), .Z(n10372) );
  MUX2_X2 U14992 ( .A(n10372), .B(n10371), .S(n10916), .Z(n10373) );
  MUX2_X2 U14993 ( .A(decode_regfile_fpregs_10__19_), .B(
        decode_regfile_fpregs_11__19_), .S(n10852), .Z(n10374) );
  MUX2_X2 U14994 ( .A(decode_regfile_fpregs_8__19_), .B(
        decode_regfile_fpregs_9__19_), .S(n10852), .Z(n10375) );
  MUX2_X2 U14995 ( .A(n10375), .B(n10374), .S(n10917), .Z(n10376) );
  MUX2_X2 U14996 ( .A(n10376), .B(n10373), .S(n10940), .Z(n10377) );
  MUX2_X2 U14997 ( .A(decode_regfile_fpregs_6__19_), .B(
        decode_regfile_fpregs_7__19_), .S(n10852), .Z(n10378) );
  MUX2_X2 U14998 ( .A(decode_regfile_fpregs_4__19_), .B(
        decode_regfile_fpregs_5__19_), .S(n10852), .Z(n10379) );
  MUX2_X2 U14999 ( .A(n10379), .B(n10378), .S(n10917), .Z(n10380) );
  MUX2_X2 U15000 ( .A(decode_regfile_fpregs_2__19_), .B(
        decode_regfile_fpregs_3__19_), .S(n10852), .Z(n10381) );
  MUX2_X2 U15001 ( .A(decode_regfile_fpregs_0__19_), .B(
        decode_regfile_fpregs_1__19_), .S(n10852), .Z(n10382) );
  MUX2_X2 U15002 ( .A(n10382), .B(n10381), .S(n10917), .Z(n10383) );
  MUX2_X2 U15003 ( .A(n10383), .B(n10380), .S(n10940), .Z(n10384) );
  MUX2_X2 U15004 ( .A(n10384), .B(n10377), .S(n10952), .Z(n10385) );
  MUX2_X2 U15005 ( .A(n10385), .B(n10370), .S(n10959), .Z(decode_regfile_N40)
         );
  MUX2_X2 U15006 ( .A(decode_regfile_fpregs_30__20_), .B(
        decode_regfile_fpregs_31__20_), .S(n10852), .Z(n10386) );
  MUX2_X2 U15007 ( .A(decode_regfile_fpregs_28__20_), .B(
        decode_regfile_fpregs_29__20_), .S(n10852), .Z(n10387) );
  MUX2_X2 U15008 ( .A(n10387), .B(n10386), .S(n10917), .Z(n10388) );
  MUX2_X2 U15009 ( .A(decode_regfile_fpregs_26__20_), .B(
        decode_regfile_fpregs_27__20_), .S(n10852), .Z(n10389) );
  MUX2_X2 U15010 ( .A(decode_regfile_fpregs_24__20_), .B(
        decode_regfile_fpregs_25__20_), .S(n10852), .Z(n10390) );
  MUX2_X2 U15011 ( .A(n10390), .B(n10389), .S(n10917), .Z(n10391) );
  MUX2_X2 U15012 ( .A(n10391), .B(n10388), .S(n10940), .Z(n10392) );
  MUX2_X2 U15013 ( .A(decode_regfile_fpregs_22__20_), .B(
        decode_regfile_fpregs_23__20_), .S(n10852), .Z(n10393) );
  MUX2_X2 U15014 ( .A(decode_regfile_fpregs_20__20_), .B(
        decode_regfile_fpregs_21__20_), .S(n10853), .Z(n10394) );
  MUX2_X2 U15015 ( .A(n10394), .B(n10393), .S(n10917), .Z(n10395) );
  MUX2_X2 U15016 ( .A(decode_regfile_fpregs_18__20_), .B(
        decode_regfile_fpregs_19__20_), .S(n10853), .Z(n10396) );
  MUX2_X2 U15017 ( .A(decode_regfile_fpregs_16__20_), .B(
        decode_regfile_fpregs_17__20_), .S(n10853), .Z(n10397) );
  MUX2_X2 U15018 ( .A(n10397), .B(n10396), .S(n10917), .Z(n10398) );
  MUX2_X2 U15019 ( .A(n10398), .B(n10395), .S(n10940), .Z(n10399) );
  MUX2_X2 U15020 ( .A(n10399), .B(n10392), .S(n10952), .Z(n10400) );
  MUX2_X2 U15021 ( .A(decode_regfile_fpregs_14__20_), .B(
        decode_regfile_fpregs_15__20_), .S(n10853), .Z(n10401) );
  MUX2_X2 U15022 ( .A(decode_regfile_fpregs_12__20_), .B(
        decode_regfile_fpregs_13__20_), .S(n10853), .Z(n10402) );
  MUX2_X2 U15023 ( .A(n10402), .B(n10401), .S(n10917), .Z(n10403) );
  MUX2_X2 U15024 ( .A(decode_regfile_fpregs_10__20_), .B(
        decode_regfile_fpregs_11__20_), .S(n10853), .Z(n10404) );
  MUX2_X2 U15025 ( .A(decode_regfile_fpregs_8__20_), .B(
        decode_regfile_fpregs_9__20_), .S(n10853), .Z(n10405) );
  MUX2_X2 U15026 ( .A(n10405), .B(n10404), .S(n10917), .Z(n10406) );
  MUX2_X2 U15027 ( .A(n10406), .B(n10403), .S(n10940), .Z(n10407) );
  MUX2_X2 U15028 ( .A(decode_regfile_fpregs_6__20_), .B(
        decode_regfile_fpregs_7__20_), .S(n10853), .Z(n10408) );
  MUX2_X2 U15029 ( .A(decode_regfile_fpregs_4__20_), .B(
        decode_regfile_fpregs_5__20_), .S(n10853), .Z(n10409) );
  MUX2_X2 U15030 ( .A(n10409), .B(n10408), .S(n10917), .Z(n10410) );
  MUX2_X2 U15031 ( .A(decode_regfile_fpregs_2__20_), .B(
        decode_regfile_fpregs_3__20_), .S(n10853), .Z(n10411) );
  MUX2_X2 U15032 ( .A(decode_regfile_fpregs_0__20_), .B(
        decode_regfile_fpregs_1__20_), .S(n10853), .Z(n10412) );
  MUX2_X2 U15033 ( .A(n10412), .B(n10411), .S(n10917), .Z(n10413) );
  MUX2_X2 U15034 ( .A(n10413), .B(n10410), .S(n10940), .Z(n10414) );
  MUX2_X2 U15035 ( .A(n10414), .B(n10407), .S(n10952), .Z(n10415) );
  MUX2_X2 U15036 ( .A(n10415), .B(n10400), .S(n10959), .Z(decode_regfile_N39)
         );
  MUX2_X2 U15037 ( .A(decode_regfile_fpregs_30__21_), .B(
        decode_regfile_fpregs_31__21_), .S(n10854), .Z(n10416) );
  MUX2_X2 U15038 ( .A(decode_regfile_fpregs_28__21_), .B(
        decode_regfile_fpregs_29__21_), .S(n10854), .Z(n10417) );
  MUX2_X2 U15039 ( .A(n10417), .B(n10416), .S(n10918), .Z(n10418) );
  MUX2_X2 U15040 ( .A(decode_regfile_fpregs_26__21_), .B(
        decode_regfile_fpregs_27__21_), .S(n10854), .Z(n10419) );
  MUX2_X2 U15041 ( .A(decode_regfile_fpregs_24__21_), .B(
        decode_regfile_fpregs_25__21_), .S(n10854), .Z(n10420) );
  MUX2_X2 U15042 ( .A(n10420), .B(n10419), .S(n10918), .Z(n10421) );
  MUX2_X2 U15043 ( .A(n10421), .B(n10418), .S(n10941), .Z(n10422) );
  MUX2_X2 U15044 ( .A(decode_regfile_fpregs_22__21_), .B(
        decode_regfile_fpregs_23__21_), .S(n10854), .Z(n10423) );
  MUX2_X2 U15045 ( .A(decode_regfile_fpregs_20__21_), .B(
        decode_regfile_fpregs_21__21_), .S(n10854), .Z(n10424) );
  MUX2_X2 U15046 ( .A(n10424), .B(n10423), .S(n10918), .Z(n10425) );
  MUX2_X2 U15047 ( .A(decode_regfile_fpregs_18__21_), .B(
        decode_regfile_fpregs_19__21_), .S(n10854), .Z(n10426) );
  MUX2_X2 U15048 ( .A(decode_regfile_fpregs_16__21_), .B(
        decode_regfile_fpregs_17__21_), .S(n10854), .Z(n10427) );
  MUX2_X2 U15049 ( .A(n10427), .B(n10426), .S(n10918), .Z(n10428) );
  MUX2_X2 U15050 ( .A(n10428), .B(n10425), .S(n10941), .Z(n10429) );
  MUX2_X2 U15051 ( .A(n10429), .B(n10422), .S(n10953), .Z(n10430) );
  MUX2_X2 U15052 ( .A(decode_regfile_fpregs_14__21_), .B(
        decode_regfile_fpregs_15__21_), .S(n10854), .Z(n10431) );
  MUX2_X2 U15053 ( .A(decode_regfile_fpregs_12__21_), .B(
        decode_regfile_fpregs_13__21_), .S(n10854), .Z(n10432) );
  MUX2_X2 U15054 ( .A(n10432), .B(n10431), .S(n10918), .Z(n10433) );
  MUX2_X2 U15055 ( .A(decode_regfile_fpregs_10__21_), .B(
        decode_regfile_fpregs_11__21_), .S(n10854), .Z(n10434) );
  MUX2_X2 U15056 ( .A(decode_regfile_fpregs_8__21_), .B(
        decode_regfile_fpregs_9__21_), .S(n10855), .Z(n10435) );
  MUX2_X2 U15057 ( .A(n10435), .B(n10434), .S(n10918), .Z(n10436) );
  MUX2_X2 U15058 ( .A(n10436), .B(n10433), .S(n10941), .Z(n10437) );
  MUX2_X2 U15059 ( .A(decode_regfile_fpregs_6__21_), .B(
        decode_regfile_fpregs_7__21_), .S(n10855), .Z(n10438) );
  MUX2_X2 U15060 ( .A(decode_regfile_fpregs_4__21_), .B(
        decode_regfile_fpregs_5__21_), .S(n10855), .Z(n10439) );
  MUX2_X2 U15061 ( .A(n10439), .B(n10438), .S(n10918), .Z(n10440) );
  MUX2_X2 U15062 ( .A(decode_regfile_fpregs_2__21_), .B(
        decode_regfile_fpregs_3__21_), .S(n10855), .Z(n10441) );
  MUX2_X2 U15063 ( .A(decode_regfile_fpregs_0__21_), .B(
        decode_regfile_fpregs_1__21_), .S(n10855), .Z(n10442) );
  MUX2_X2 U15064 ( .A(n10442), .B(n10441), .S(n10918), .Z(n10443) );
  MUX2_X2 U15065 ( .A(n10443), .B(n10440), .S(n10941), .Z(n10444) );
  MUX2_X2 U15066 ( .A(n10444), .B(n10437), .S(n10953), .Z(n10445) );
  MUX2_X2 U15067 ( .A(n10445), .B(n10430), .S(n10960), .Z(decode_regfile_N38)
         );
  MUX2_X2 U15068 ( .A(decode_regfile_fpregs_30__22_), .B(
        decode_regfile_fpregs_31__22_), .S(n10855), .Z(n10446) );
  MUX2_X2 U15069 ( .A(decode_regfile_fpregs_28__22_), .B(
        decode_regfile_fpregs_29__22_), .S(n10855), .Z(n10447) );
  MUX2_X2 U15070 ( .A(n10447), .B(n10446), .S(n10918), .Z(n10448) );
  MUX2_X2 U15071 ( .A(decode_regfile_fpregs_26__22_), .B(
        decode_regfile_fpregs_27__22_), .S(n10855), .Z(n10449) );
  MUX2_X2 U15072 ( .A(decode_regfile_fpregs_24__22_), .B(
        decode_regfile_fpregs_25__22_), .S(n10855), .Z(n10450) );
  MUX2_X2 U15073 ( .A(n10450), .B(n10449), .S(n10918), .Z(n10451) );
  MUX2_X2 U15074 ( .A(n10451), .B(n10448), .S(n10941), .Z(n10452) );
  MUX2_X2 U15075 ( .A(decode_regfile_fpregs_22__22_), .B(
        decode_regfile_fpregs_23__22_), .S(n10855), .Z(n10453) );
  MUX2_X2 U15076 ( .A(decode_regfile_fpregs_20__22_), .B(
        decode_regfile_fpregs_21__22_), .S(n10855), .Z(n10454) );
  MUX2_X2 U15077 ( .A(n10454), .B(n10453), .S(n10918), .Z(n10455) );
  MUX2_X2 U15078 ( .A(decode_regfile_fpregs_18__22_), .B(
        decode_regfile_fpregs_19__22_), .S(n10856), .Z(n10456) );
  MUX2_X2 U15079 ( .A(decode_regfile_fpregs_16__22_), .B(
        decode_regfile_fpregs_17__22_), .S(n10856), .Z(n10457) );
  MUX2_X2 U15080 ( .A(n10457), .B(n10456), .S(n10919), .Z(n10458) );
  MUX2_X2 U15081 ( .A(n10458), .B(n10455), .S(n10941), .Z(n10459) );
  MUX2_X2 U15082 ( .A(n10459), .B(n10452), .S(n10953), .Z(n10460) );
  MUX2_X2 U15083 ( .A(decode_regfile_fpregs_14__22_), .B(
        decode_regfile_fpregs_15__22_), .S(n10856), .Z(n10461) );
  MUX2_X2 U15084 ( .A(decode_regfile_fpregs_12__22_), .B(
        decode_regfile_fpregs_13__22_), .S(n10856), .Z(n10462) );
  MUX2_X2 U15085 ( .A(n10462), .B(n10461), .S(n10919), .Z(n10463) );
  MUX2_X2 U15086 ( .A(decode_regfile_fpregs_10__22_), .B(
        decode_regfile_fpregs_11__22_), .S(n10856), .Z(n10464) );
  MUX2_X2 U15087 ( .A(decode_regfile_fpregs_8__22_), .B(
        decode_regfile_fpregs_9__22_), .S(n10856), .Z(n10465) );
  MUX2_X2 U15088 ( .A(n10465), .B(n10464), .S(n10919), .Z(n10466) );
  MUX2_X2 U15089 ( .A(n10466), .B(n10463), .S(n10941), .Z(n10467) );
  MUX2_X2 U15090 ( .A(decode_regfile_fpregs_6__22_), .B(
        decode_regfile_fpregs_7__22_), .S(n10856), .Z(n10468) );
  MUX2_X2 U15091 ( .A(decode_regfile_fpregs_4__22_), .B(
        decode_regfile_fpregs_5__22_), .S(n10856), .Z(n10469) );
  MUX2_X2 U15092 ( .A(n10469), .B(n10468), .S(n10919), .Z(n10470) );
  MUX2_X2 U15093 ( .A(decode_regfile_fpregs_2__22_), .B(
        decode_regfile_fpregs_3__22_), .S(n10856), .Z(n10471) );
  MUX2_X2 U15094 ( .A(decode_regfile_fpregs_0__22_), .B(
        decode_regfile_fpregs_1__22_), .S(n10856), .Z(n10472) );
  MUX2_X2 U15095 ( .A(n10472), .B(n10471), .S(n10919), .Z(n10473) );
  MUX2_X2 U15096 ( .A(n10473), .B(n10470), .S(n10941), .Z(n10474) );
  MUX2_X2 U15097 ( .A(n10474), .B(n10467), .S(n10953), .Z(n10475) );
  MUX2_X2 U15098 ( .A(n10475), .B(n10460), .S(n10960), .Z(decode_regfile_N37)
         );
  MUX2_X2 U15099 ( .A(decode_regfile_fpregs_30__23_), .B(
        decode_regfile_fpregs_31__23_), .S(n10856), .Z(n10476) );
  MUX2_X2 U15100 ( .A(decode_regfile_fpregs_28__23_), .B(
        decode_regfile_fpregs_29__23_), .S(n10857), .Z(n10477) );
  MUX2_X2 U15101 ( .A(n10477), .B(n10476), .S(n10919), .Z(n10478) );
  MUX2_X2 U15102 ( .A(decode_regfile_fpregs_26__23_), .B(
        decode_regfile_fpregs_27__23_), .S(n10857), .Z(n10479) );
  MUX2_X2 U15103 ( .A(decode_regfile_fpregs_24__23_), .B(
        decode_regfile_fpregs_25__23_), .S(n10857), .Z(n10480) );
  MUX2_X2 U15104 ( .A(n10480), .B(n10479), .S(n10919), .Z(n10481) );
  MUX2_X2 U15105 ( .A(n10481), .B(n10478), .S(n10941), .Z(n10482) );
  MUX2_X2 U15106 ( .A(decode_regfile_fpregs_22__23_), .B(
        decode_regfile_fpregs_23__23_), .S(n10857), .Z(n10483) );
  MUX2_X2 U15107 ( .A(decode_regfile_fpregs_20__23_), .B(
        decode_regfile_fpregs_21__23_), .S(n10857), .Z(n10484) );
  MUX2_X2 U15108 ( .A(n10484), .B(n10483), .S(n10919), .Z(n10485) );
  MUX2_X2 U15109 ( .A(decode_regfile_fpregs_18__23_), .B(
        decode_regfile_fpregs_19__23_), .S(n10857), .Z(n10486) );
  MUX2_X2 U15110 ( .A(decode_regfile_fpregs_16__23_), .B(
        decode_regfile_fpregs_17__23_), .S(n10857), .Z(n10487) );
  MUX2_X2 U15111 ( .A(n10487), .B(n10486), .S(n10919), .Z(n10488) );
  MUX2_X2 U15112 ( .A(n10488), .B(n10485), .S(n10941), .Z(n10489) );
  MUX2_X2 U15113 ( .A(n10489), .B(n10482), .S(n10953), .Z(n10490) );
  MUX2_X2 U15114 ( .A(decode_regfile_fpregs_14__23_), .B(
        decode_regfile_fpregs_15__23_), .S(n10857), .Z(n10491) );
  MUX2_X2 U15115 ( .A(decode_regfile_fpregs_12__23_), .B(
        decode_regfile_fpregs_13__23_), .S(n10857), .Z(n10492) );
  MUX2_X2 U15116 ( .A(n10492), .B(n10491), .S(n10919), .Z(n10493) );
  MUX2_X2 U15117 ( .A(decode_regfile_fpregs_10__23_), .B(
        decode_regfile_fpregs_11__23_), .S(n10857), .Z(n10494) );
  MUX2_X2 U15118 ( .A(decode_regfile_fpregs_8__23_), .B(
        decode_regfile_fpregs_9__23_), .S(n10857), .Z(n10495) );
  MUX2_X2 U15119 ( .A(n10495), .B(n10494), .S(n10919), .Z(n10496) );
  MUX2_X2 U15120 ( .A(n10496), .B(n10493), .S(n10941), .Z(n10497) );
  MUX2_X2 U15121 ( .A(decode_regfile_fpregs_6__23_), .B(
        decode_regfile_fpregs_7__23_), .S(n10858), .Z(n10498) );
  MUX2_X2 U15122 ( .A(decode_regfile_fpregs_4__23_), .B(
        decode_regfile_fpregs_5__23_), .S(n10858), .Z(n10499) );
  MUX2_X2 U15123 ( .A(n10499), .B(n10498), .S(n10870), .Z(n10500) );
  MUX2_X2 U15124 ( .A(decode_regfile_fpregs_2__23_), .B(
        decode_regfile_fpregs_3__23_), .S(n10858), .Z(n10501) );
  MUX2_X2 U15125 ( .A(decode_regfile_fpregs_0__23_), .B(
        decode_regfile_fpregs_1__23_), .S(n10858), .Z(n10502) );
  MUX2_X2 U15126 ( .A(n10502), .B(n10501), .S(n10864), .Z(n10503) );
  MUX2_X2 U15127 ( .A(n10503), .B(n10500), .S(n10942), .Z(n10504) );
  MUX2_X2 U15128 ( .A(n10504), .B(n10497), .S(n10953), .Z(n10505) );
  MUX2_X2 U15129 ( .A(n10505), .B(n10490), .S(n10960), .Z(decode_regfile_N36)
         );
  MUX2_X2 U15130 ( .A(decode_regfile_fpregs_30__24_), .B(
        decode_regfile_fpregs_31__24_), .S(n10858), .Z(n10506) );
  MUX2_X2 U15131 ( .A(decode_regfile_fpregs_28__24_), .B(
        decode_regfile_fpregs_29__24_), .S(n10858), .Z(n10507) );
  MUX2_X2 U15132 ( .A(n10507), .B(n10506), .S(n10865), .Z(n10508) );
  MUX2_X2 U15133 ( .A(decode_regfile_fpregs_26__24_), .B(
        decode_regfile_fpregs_27__24_), .S(n10858), .Z(n10509) );
  MUX2_X2 U15134 ( .A(decode_regfile_fpregs_24__24_), .B(
        decode_regfile_fpregs_25__24_), .S(n10858), .Z(n10510) );
  MUX2_X2 U15135 ( .A(n10510), .B(n10509), .S(n10868), .Z(n10511) );
  MUX2_X2 U15136 ( .A(n10511), .B(n10508), .S(n10942), .Z(n10512) );
  MUX2_X2 U15137 ( .A(decode_regfile_fpregs_22__24_), .B(
        decode_regfile_fpregs_23__24_), .S(n10858), .Z(n10513) );
  MUX2_X2 U15138 ( .A(decode_regfile_fpregs_20__24_), .B(
        decode_regfile_fpregs_21__24_), .S(n10858), .Z(n10514) );
  MUX2_X2 U15139 ( .A(n10514), .B(n10513), .S(n10869), .Z(n10515) );
  MUX2_X2 U15140 ( .A(decode_regfile_fpregs_18__24_), .B(
        decode_regfile_fpregs_19__24_), .S(n10858), .Z(n10516) );
  MUX2_X2 U15141 ( .A(decode_regfile_fpregs_16__24_), .B(
        decode_regfile_fpregs_17__24_), .S(n10756), .Z(n10517) );
  MUX2_X2 U15142 ( .A(n10517), .B(n10516), .S(n10863), .Z(n10518) );
  MUX2_X2 U15143 ( .A(n10518), .B(n10515), .S(n10942), .Z(n10519) );
  MUX2_X2 U15144 ( .A(n10519), .B(n10512), .S(n10953), .Z(n10520) );
  MUX2_X2 U15145 ( .A(decode_regfile_fpregs_14__24_), .B(
        decode_regfile_fpregs_15__24_), .S(n10758), .Z(n10521) );
  MUX2_X2 U15146 ( .A(decode_regfile_fpregs_12__24_), .B(
        decode_regfile_fpregs_13__24_), .S(n10759), .Z(n10522) );
  MUX2_X2 U15147 ( .A(n10522), .B(n10521), .S(n10867), .Z(n10523) );
  MUX2_X2 U15148 ( .A(decode_regfile_fpregs_10__24_), .B(
        decode_regfile_fpregs_11__24_), .S(n10754), .Z(n10524) );
  MUX2_X2 U15149 ( .A(decode_regfile_fpregs_8__24_), .B(
        decode_regfile_fpregs_9__24_), .S(n10760), .Z(n10525) );
  MUX2_X2 U15150 ( .A(n10525), .B(n10524), .S(n10865), .Z(n10526) );
  MUX2_X2 U15151 ( .A(n10526), .B(n10523), .S(n10942), .Z(n10527) );
  MUX2_X2 U15152 ( .A(decode_regfile_fpregs_6__24_), .B(
        decode_regfile_fpregs_7__24_), .S(n10753), .Z(n10528) );
  MUX2_X2 U15153 ( .A(decode_regfile_fpregs_4__24_), .B(
        decode_regfile_fpregs_5__24_), .S(n10755), .Z(n10529) );
  MUX2_X2 U15154 ( .A(n10529), .B(n10528), .S(n10866), .Z(n10530) );
  MUX2_X2 U15155 ( .A(decode_regfile_fpregs_2__24_), .B(
        decode_regfile_fpregs_3__24_), .S(n10751), .Z(n10531) );
  MUX2_X2 U15156 ( .A(decode_regfile_fpregs_0__24_), .B(
        decode_regfile_fpregs_1__24_), .S(n10752), .Z(n10532) );
  MUX2_X2 U15157 ( .A(n10532), .B(n10531), .S(n10873), .Z(n10533) );
  MUX2_X2 U15158 ( .A(n10533), .B(n10530), .S(n10942), .Z(n10534) );
  MUX2_X2 U15159 ( .A(n10534), .B(n10527), .S(n10953), .Z(n10535) );
  MUX2_X2 U15160 ( .A(n10535), .B(n10520), .S(n10960), .Z(decode_regfile_N35)
         );
  MUX2_X2 U15161 ( .A(decode_regfile_fpregs_30__25_), .B(
        decode_regfile_fpregs_31__25_), .S(n10749), .Z(n10536) );
  MUX2_X2 U15162 ( .A(decode_regfile_fpregs_28__25_), .B(
        decode_regfile_fpregs_29__25_), .S(n10750), .Z(n10537) );
  MUX2_X2 U15163 ( .A(n10537), .B(n10536), .S(n10874), .Z(n10538) );
  MUX2_X2 U15164 ( .A(decode_regfile_fpregs_26__25_), .B(
        decode_regfile_fpregs_27__25_), .S(n10859), .Z(n10539) );
  MUX2_X2 U15165 ( .A(decode_regfile_fpregs_24__25_), .B(
        decode_regfile_fpregs_25__25_), .S(n10859), .Z(n10540) );
  MUX2_X2 U15166 ( .A(n10540), .B(n10539), .S(n10920), .Z(n10541) );
  MUX2_X2 U15167 ( .A(n10541), .B(n10538), .S(n10942), .Z(n10542) );
  MUX2_X2 U15168 ( .A(decode_regfile_fpregs_22__25_), .B(
        decode_regfile_fpregs_23__25_), .S(n10859), .Z(n10543) );
  MUX2_X2 U15169 ( .A(decode_regfile_fpregs_20__25_), .B(
        decode_regfile_fpregs_21__25_), .S(n10859), .Z(n10544) );
  MUX2_X2 U15170 ( .A(n10544), .B(n10543), .S(n10920), .Z(n10545) );
  MUX2_X2 U15171 ( .A(decode_regfile_fpregs_18__25_), .B(
        decode_regfile_fpregs_19__25_), .S(n10859), .Z(n10546) );
  MUX2_X2 U15172 ( .A(decode_regfile_fpregs_16__25_), .B(
        decode_regfile_fpregs_17__25_), .S(n10859), .Z(n10547) );
  MUX2_X2 U15173 ( .A(n10547), .B(n10546), .S(n10920), .Z(n10548) );
  MUX2_X2 U15174 ( .A(n10548), .B(n10545), .S(n10942), .Z(n10549) );
  MUX2_X2 U15175 ( .A(n10549), .B(n10542), .S(n10953), .Z(n10550) );
  MUX2_X2 U15176 ( .A(decode_regfile_fpregs_14__25_), .B(
        decode_regfile_fpregs_15__25_), .S(n10859), .Z(n10551) );
  MUX2_X2 U15177 ( .A(decode_regfile_fpregs_12__25_), .B(
        decode_regfile_fpregs_13__25_), .S(n10859), .Z(n10552) );
  MUX2_X2 U15178 ( .A(n10552), .B(n10551), .S(n10920), .Z(n10553) );
  MUX2_X2 U15179 ( .A(decode_regfile_fpregs_10__25_), .B(
        decode_regfile_fpregs_11__25_), .S(n10859), .Z(n10554) );
  MUX2_X2 U15180 ( .A(decode_regfile_fpregs_8__25_), .B(
        decode_regfile_fpregs_9__25_), .S(n10859), .Z(n10555) );
  MUX2_X2 U15181 ( .A(n10555), .B(n10554), .S(n10920), .Z(n10556) );
  MUX2_X2 U15182 ( .A(n10556), .B(n10553), .S(n10942), .Z(n10557) );
  MUX2_X2 U15183 ( .A(decode_regfile_fpregs_6__25_), .B(
        decode_regfile_fpregs_7__25_), .S(n10859), .Z(n10558) );
  MUX2_X2 U15184 ( .A(decode_regfile_fpregs_4__25_), .B(
        decode_regfile_fpregs_5__25_), .S(n10860), .Z(n10559) );
  MUX2_X2 U15185 ( .A(n10559), .B(n10558), .S(n10920), .Z(n10560) );
  MUX2_X2 U15186 ( .A(decode_regfile_fpregs_2__25_), .B(
        decode_regfile_fpregs_3__25_), .S(n10860), .Z(n10561) );
  MUX2_X2 U15187 ( .A(decode_regfile_fpregs_0__25_), .B(
        decode_regfile_fpregs_1__25_), .S(n10860), .Z(n10562) );
  MUX2_X2 U15188 ( .A(n10562), .B(n10561), .S(n10920), .Z(n10563) );
  MUX2_X2 U15189 ( .A(n10563), .B(n10560), .S(n10942), .Z(n10564) );
  MUX2_X2 U15190 ( .A(n10564), .B(n10557), .S(n10953), .Z(n10565) );
  MUX2_X2 U15191 ( .A(n10565), .B(n10550), .S(n10960), .Z(decode_regfile_N34)
         );
  MUX2_X2 U15192 ( .A(decode_regfile_fpregs_30__26_), .B(
        decode_regfile_fpregs_31__26_), .S(n10860), .Z(n10566) );
  MUX2_X2 U15193 ( .A(decode_regfile_fpregs_28__26_), .B(
        decode_regfile_fpregs_29__26_), .S(n10860), .Z(n10567) );
  MUX2_X2 U15194 ( .A(n10567), .B(n10566), .S(n10920), .Z(n10568) );
  MUX2_X2 U15195 ( .A(decode_regfile_fpregs_26__26_), .B(
        decode_regfile_fpregs_27__26_), .S(n10860), .Z(n10569) );
  MUX2_X2 U15196 ( .A(decode_regfile_fpregs_24__26_), .B(
        decode_regfile_fpregs_25__26_), .S(n10860), .Z(n10570) );
  MUX2_X2 U15197 ( .A(n10570), .B(n10569), .S(n10920), .Z(n10571) );
  MUX2_X2 U15198 ( .A(n10571), .B(n10568), .S(n10942), .Z(n10572) );
  MUX2_X2 U15199 ( .A(decode_regfile_fpregs_22__26_), .B(
        decode_regfile_fpregs_23__26_), .S(n10860), .Z(n10573) );
  MUX2_X2 U15200 ( .A(decode_regfile_fpregs_20__26_), .B(
        decode_regfile_fpregs_21__26_), .S(n10860), .Z(n10574) );
  MUX2_X2 U15201 ( .A(n10574), .B(n10573), .S(n10920), .Z(n10575) );
  MUX2_X2 U15202 ( .A(decode_regfile_fpregs_18__26_), .B(
        decode_regfile_fpregs_19__26_), .S(n10860), .Z(n10576) );
  MUX2_X2 U15203 ( .A(decode_regfile_fpregs_16__26_), .B(
        decode_regfile_fpregs_17__26_), .S(n10860), .Z(n10577) );
  MUX2_X2 U15204 ( .A(n10577), .B(n10576), .S(n10920), .Z(n10578) );
  MUX2_X2 U15205 ( .A(n10578), .B(n10575), .S(n10942), .Z(n10579) );
  MUX2_X2 U15206 ( .A(n10579), .B(n10572), .S(n10953), .Z(n10580) );
  MUX2_X2 U15207 ( .A(decode_regfile_fpregs_14__26_), .B(
        decode_regfile_fpregs_15__26_), .S(n10861), .Z(n10581) );
  MUX2_X2 U15208 ( .A(decode_regfile_fpregs_12__26_), .B(
        decode_regfile_fpregs_13__26_), .S(n10861), .Z(n10582) );
  MUX2_X2 U15209 ( .A(n10582), .B(n10581), .S(n10866), .Z(n10583) );
  MUX2_X2 U15210 ( .A(decode_regfile_fpregs_10__26_), .B(
        decode_regfile_fpregs_11__26_), .S(n10861), .Z(n10584) );
  MUX2_X2 U15211 ( .A(decode_regfile_fpregs_8__26_), .B(
        decode_regfile_fpregs_9__26_), .S(n10861), .Z(n10585) );
  MUX2_X2 U15212 ( .A(n10585), .B(n10584), .S(n10876), .Z(n10586) );
  MUX2_X2 U15213 ( .A(n10586), .B(n10583), .S(n10921), .Z(n10587) );
  MUX2_X2 U15214 ( .A(decode_regfile_fpregs_6__26_), .B(
        decode_regfile_fpregs_7__26_), .S(n10861), .Z(n10588) );
  MUX2_X2 U15215 ( .A(decode_regfile_fpregs_4__26_), .B(
        decode_regfile_fpregs_5__26_), .S(n10861), .Z(n10589) );
  MUX2_X2 U15216 ( .A(n10589), .B(n10588), .S(n10877), .Z(n10590) );
  MUX2_X2 U15217 ( .A(decode_regfile_fpregs_2__26_), .B(
        decode_regfile_fpregs_3__26_), .S(n10861), .Z(n10591) );
  MUX2_X2 U15218 ( .A(decode_regfile_fpregs_0__26_), .B(
        decode_regfile_fpregs_1__26_), .S(n10861), .Z(n10592) );
  MUX2_X2 U15219 ( .A(n10592), .B(n10591), .S(n10871), .Z(n10593) );
  MUX2_X2 U15220 ( .A(n10593), .B(n10590), .S(n10930), .Z(n10594) );
  MUX2_X2 U15221 ( .A(n10594), .B(n10587), .S(n10954), .Z(n10595) );
  MUX2_X2 U15222 ( .A(n10595), .B(n10580), .S(n10960), .Z(decode_regfile_N33)
         );
  MUX2_X2 U15223 ( .A(decode_regfile_fpregs_30__27_), .B(
        decode_regfile_fpregs_31__27_), .S(n10861), .Z(n10596) );
  MUX2_X2 U15224 ( .A(decode_regfile_fpregs_28__27_), .B(
        decode_regfile_fpregs_29__27_), .S(n10861), .Z(n10597) );
  MUX2_X2 U15225 ( .A(n10597), .B(n10596), .S(n10864), .Z(n10598) );
  MUX2_X2 U15226 ( .A(decode_regfile_fpregs_26__27_), .B(
        decode_regfile_fpregs_27__27_), .S(n10861), .Z(n10599) );
  MUX2_X2 U15227 ( .A(decode_regfile_fpregs_24__27_), .B(
        decode_regfile_fpregs_25__27_), .S(n10754), .Z(n10600) );
  MUX2_X2 U15228 ( .A(n10600), .B(n10599), .S(n10873), .Z(n10601) );
  MUX2_X2 U15229 ( .A(n10601), .B(n10598), .S(decode_rs2_2_), .Z(n10602) );
  MUX2_X2 U15230 ( .A(decode_regfile_fpregs_22__27_), .B(
        decode_regfile_fpregs_23__27_), .S(n10747), .Z(n10603) );
  MUX2_X2 U15231 ( .A(decode_regfile_fpregs_20__27_), .B(
        decode_regfile_fpregs_21__27_), .S(n10759), .Z(n10604) );
  MUX2_X2 U15232 ( .A(n10604), .B(n10603), .S(n10863), .Z(n10605) );
  MUX2_X2 U15233 ( .A(decode_regfile_fpregs_18__27_), .B(
        decode_regfile_fpregs_19__27_), .S(n10756), .Z(n10606) );
  MUX2_X2 U15234 ( .A(decode_regfile_fpregs_16__27_), .B(
        decode_regfile_fpregs_17__27_), .S(n10752), .Z(n10607) );
  MUX2_X2 U15235 ( .A(n10607), .B(n10606), .S(n10872), .Z(n10608) );
  MUX2_X2 U15236 ( .A(n10608), .B(n10605), .S(decode_rs2_2_), .Z(n10609) );
  MUX2_X2 U15237 ( .A(n10609), .B(n10602), .S(n10954), .Z(n10610) );
  MUX2_X2 U15238 ( .A(decode_regfile_fpregs_14__27_), .B(
        decode_regfile_fpregs_15__27_), .S(n10758), .Z(n10611) );
  MUX2_X2 U15239 ( .A(decode_regfile_fpregs_12__27_), .B(
        decode_regfile_fpregs_13__27_), .S(n10753), .Z(n10612) );
  MUX2_X2 U15240 ( .A(n10612), .B(n10611), .S(n10864), .Z(n10613) );
  MUX2_X2 U15241 ( .A(decode_regfile_fpregs_10__27_), .B(
        decode_regfile_fpregs_11__27_), .S(n10760), .Z(n10614) );
  MUX2_X2 U15242 ( .A(decode_regfile_fpregs_8__27_), .B(
        decode_regfile_fpregs_9__27_), .S(n10776), .Z(n10615) );
  MUX2_X2 U15243 ( .A(n10615), .B(n10614), .S(n10878), .Z(n10616) );
  MUX2_X2 U15244 ( .A(n10616), .B(n10613), .S(n10921), .Z(n10617) );
  MUX2_X2 U15245 ( .A(decode_regfile_fpregs_6__27_), .B(
        decode_regfile_fpregs_7__27_), .S(n10755), .Z(n10618) );
  MUX2_X2 U15246 ( .A(decode_regfile_fpregs_4__27_), .B(
        decode_regfile_fpregs_5__27_), .S(n10751), .Z(n10619) );
  MUX2_X2 U15247 ( .A(n10619), .B(n10618), .S(n10875), .Z(n10620) );
  MUX2_X2 U15248 ( .A(decode_regfile_fpregs_2__27_), .B(
        decode_regfile_fpregs_3__27_), .S(n10862), .Z(n10621) );
  MUX2_X2 U15249 ( .A(decode_regfile_fpregs_0__27_), .B(
        decode_regfile_fpregs_1__27_), .S(n10862), .Z(n10622) );
  MUX2_X2 U15250 ( .A(n10622), .B(n10621), .S(n10873), .Z(n10623) );
  MUX2_X2 U15251 ( .A(n10623), .B(n10620), .S(n10929), .Z(n10624) );
  MUX2_X2 U15252 ( .A(n10624), .B(n10617), .S(n10954), .Z(n10625) );
  MUX2_X2 U15253 ( .A(n10625), .B(n10610), .S(n10960), .Z(decode_regfile_N32)
         );
  MUX2_X2 U15254 ( .A(decode_regfile_fpregs_30__28_), .B(
        decode_regfile_fpregs_31__28_), .S(n10862), .Z(n10626) );
  MUX2_X2 U15255 ( .A(decode_regfile_fpregs_28__28_), .B(
        decode_regfile_fpregs_29__28_), .S(n10862), .Z(n10627) );
  MUX2_X2 U15256 ( .A(n10627), .B(n10626), .S(n10864), .Z(n10628) );
  MUX2_X2 U15257 ( .A(decode_regfile_fpregs_26__28_), .B(
        decode_regfile_fpregs_27__28_), .S(n10862), .Z(n10629) );
  MUX2_X2 U15258 ( .A(decode_regfile_fpregs_24__28_), .B(
        decode_regfile_fpregs_25__28_), .S(n10862), .Z(n10630) );
  MUX2_X2 U15259 ( .A(n10630), .B(n10629), .S(n10868), .Z(n10631) );
  MUX2_X2 U15260 ( .A(n10631), .B(n10628), .S(n10921), .Z(n10632) );
  MUX2_X2 U15261 ( .A(decode_regfile_fpregs_22__28_), .B(
        decode_regfile_fpregs_23__28_), .S(n10862), .Z(n10633) );
  MUX2_X2 U15262 ( .A(decode_regfile_fpregs_20__28_), .B(
        decode_regfile_fpregs_21__28_), .S(n10862), .Z(n10634) );
  MUX2_X2 U15263 ( .A(n10634), .B(n10633), .S(n10869), .Z(n10635) );
  MUX2_X2 U15264 ( .A(decode_regfile_fpregs_18__28_), .B(
        decode_regfile_fpregs_19__28_), .S(n10862), .Z(n10636) );
  MUX2_X2 U15265 ( .A(decode_regfile_fpregs_16__28_), .B(
        decode_regfile_fpregs_17__28_), .S(n10862), .Z(n10637) );
  MUX2_X2 U15266 ( .A(n10637), .B(n10636), .S(n10864), .Z(n10638) );
  MUX2_X2 U15267 ( .A(n10638), .B(n10635), .S(decode_rs2_2_), .Z(n10639) );
  MUX2_X2 U15268 ( .A(n10639), .B(n10632), .S(n10954), .Z(n10640) );
  MUX2_X2 U15269 ( .A(decode_regfile_fpregs_14__28_), .B(
        decode_regfile_fpregs_15__28_), .S(n10862), .Z(n10641) );
  MUX2_X2 U15270 ( .A(decode_regfile_fpregs_12__28_), .B(
        decode_regfile_fpregs_13__28_), .S(n10771), .Z(n10642) );
  MUX2_X2 U15271 ( .A(n10642), .B(n10641), .S(n10867), .Z(n10643) );
  MUX2_X2 U15272 ( .A(decode_regfile_fpregs_10__28_), .B(
        decode_regfile_fpregs_11__28_), .S(n10761), .Z(n10644) );
  MUX2_X2 U15273 ( .A(decode_regfile_fpregs_8__28_), .B(
        decode_regfile_fpregs_9__28_), .S(n10768), .Z(n10645) );
  MUX2_X2 U15274 ( .A(n10645), .B(n10644), .S(n10863), .Z(n10646) );
  MUX2_X2 U15275 ( .A(n10646), .B(n10643), .S(n10924), .Z(n10647) );
  MUX2_X2 U15276 ( .A(decode_regfile_fpregs_6__28_), .B(
        decode_regfile_fpregs_7__28_), .S(n10762), .Z(n10648) );
  MUX2_X2 U15277 ( .A(decode_regfile_fpregs_4__28_), .B(
        decode_regfile_fpregs_5__28_), .S(n10767), .Z(n10649) );
  MUX2_X2 U15278 ( .A(n10649), .B(n10648), .S(n10866), .Z(n10650) );
  MUX2_X2 U15279 ( .A(decode_regfile_fpregs_2__28_), .B(
        decode_regfile_fpregs_3__28_), .S(n10757), .Z(n10651) );
  MUX2_X2 U15280 ( .A(decode_regfile_fpregs_0__28_), .B(
        decode_regfile_fpregs_1__28_), .S(n10748), .Z(n10652) );
  MUX2_X2 U15281 ( .A(n10652), .B(n10651), .S(n10877), .Z(n10653) );
  MUX2_X2 U15282 ( .A(n10653), .B(n10650), .S(n10923), .Z(n10654) );
  MUX2_X2 U15283 ( .A(n10654), .B(n10647), .S(n10954), .Z(n10655) );
  MUX2_X2 U15284 ( .A(n10655), .B(n10640), .S(n10960), .Z(decode_regfile_N31)
         );
  MUX2_X2 U15285 ( .A(decode_regfile_fpregs_30__29_), .B(
        decode_regfile_fpregs_31__29_), .S(n10747), .Z(n10656) );
  MUX2_X2 U15286 ( .A(decode_regfile_fpregs_28__29_), .B(
        decode_regfile_fpregs_29__29_), .S(n10769), .Z(n10657) );
  MUX2_X2 U15287 ( .A(n10657), .B(n10656), .S(n10865), .Z(n10658) );
  MUX2_X2 U15288 ( .A(decode_regfile_fpregs_26__29_), .B(
        decode_regfile_fpregs_27__29_), .S(n10770), .Z(n10659) );
  MUX2_X2 U15289 ( .A(decode_regfile_fpregs_24__29_), .B(
        decode_regfile_fpregs_25__29_), .S(n10763), .Z(n10660) );
  MUX2_X2 U15290 ( .A(n10660), .B(n10659), .S(n10870), .Z(n10661) );
  MUX2_X2 U15291 ( .A(n10661), .B(n10658), .S(decode_rs2_2_), .Z(n10662) );
  MUX2_X2 U15292 ( .A(decode_regfile_fpregs_22__29_), .B(
        decode_regfile_fpregs_23__29_), .S(n10746), .Z(n10663) );
  MUX2_X2 U15293 ( .A(decode_regfile_fpregs_20__29_), .B(
        decode_regfile_fpregs_21__29_), .S(n10762), .Z(n10664) );
  MUX2_X2 U15294 ( .A(n10664), .B(n10663), .S(n10876), .Z(n10665) );
  MUX2_X2 U15295 ( .A(decode_regfile_fpregs_18__29_), .B(
        decode_regfile_fpregs_19__29_), .S(n10767), .Z(n10666) );
  MUX2_X2 U15296 ( .A(decode_regfile_fpregs_16__29_), .B(
        decode_regfile_fpregs_17__29_), .S(n10748), .Z(n10667) );
  MUX2_X2 U15297 ( .A(n10667), .B(n10666), .S(n10869), .Z(n10668) );
  MUX2_X2 U15298 ( .A(n10668), .B(n10665), .S(n10921), .Z(n10669) );
  MUX2_X2 U15299 ( .A(n10669), .B(n10662), .S(n10954), .Z(n10670) );
  MUX2_X2 U15300 ( .A(decode_regfile_fpregs_14__29_), .B(
        decode_regfile_fpregs_15__29_), .S(n10771), .Z(n10671) );
  MUX2_X2 U15301 ( .A(decode_regfile_fpregs_12__29_), .B(
        decode_regfile_fpregs_13__29_), .S(n10763), .Z(n10672) );
  MUX2_X2 U15302 ( .A(n10672), .B(n10671), .S(n10872), .Z(n10673) );
  MUX2_X2 U15303 ( .A(decode_regfile_fpregs_10__29_), .B(
        decode_regfile_fpregs_11__29_), .S(n10768), .Z(n10674) );
  MUX2_X2 U15304 ( .A(decode_regfile_fpregs_8__29_), .B(
        decode_regfile_fpregs_9__29_), .S(n10749), .Z(n10675) );
  MUX2_X2 U15305 ( .A(n10675), .B(n10674), .S(n10867), .Z(n10676) );
  MUX2_X2 U15306 ( .A(n10676), .B(n10673), .S(decode_rs2_2_), .Z(n10677) );
  MUX2_X2 U15307 ( .A(decode_regfile_fpregs_6__29_), .B(
        decode_regfile_fpregs_7__29_), .S(n10761), .Z(n10678) );
  MUX2_X2 U15308 ( .A(decode_regfile_fpregs_4__29_), .B(
        decode_regfile_fpregs_5__29_), .S(n10757), .Z(n10679) );
  MUX2_X2 U15309 ( .A(n10679), .B(n10678), .S(n10865), .Z(n10680) );
  MUX2_X2 U15310 ( .A(decode_regfile_fpregs_2__29_), .B(
        decode_regfile_fpregs_3__29_), .S(n10750), .Z(n10681) );
  MUX2_X2 U15311 ( .A(decode_regfile_fpregs_0__29_), .B(
        decode_regfile_fpregs_1__29_), .S(n10774), .Z(n10682) );
  MUX2_X2 U15312 ( .A(n10682), .B(n10681), .S(n10870), .Z(n10683) );
  MUX2_X2 U15313 ( .A(n10683), .B(n10680), .S(n10921), .Z(n10684) );
  MUX2_X2 U15314 ( .A(n10684), .B(n10677), .S(n10954), .Z(n10685) );
  MUX2_X2 U15315 ( .A(n10685), .B(n10670), .S(n10960), .Z(decode_regfile_N30)
         );
  MUX2_X2 U15316 ( .A(decode_regfile_fpregs_30__30_), .B(
        decode_regfile_fpregs_31__30_), .S(n10746), .Z(n10686) );
  MUX2_X2 U15317 ( .A(decode_regfile_fpregs_28__30_), .B(
        decode_regfile_fpregs_29__30_), .S(n10776), .Z(n10687) );
  MUX2_X2 U15318 ( .A(n10687), .B(n10686), .S(n10875), .Z(n10688) );
  MUX2_X2 U15319 ( .A(decode_regfile_fpregs_26__30_), .B(
        decode_regfile_fpregs_27__30_), .S(n10747), .Z(n10689) );
  MUX2_X2 U15320 ( .A(decode_regfile_fpregs_24__30_), .B(
        decode_regfile_fpregs_25__30_), .S(n10766), .Z(n10690) );
  MUX2_X2 U15321 ( .A(n10690), .B(n10689), .S(n10874), .Z(n10691) );
  MUX2_X2 U15322 ( .A(n10691), .B(n10688), .S(decode_rs2_2_), .Z(n10692) );
  MUX2_X2 U15323 ( .A(decode_regfile_fpregs_22__30_), .B(
        decode_regfile_fpregs_23__30_), .S(n10749), .Z(n10693) );
  MUX2_X2 U15324 ( .A(decode_regfile_fpregs_20__30_), .B(
        decode_regfile_fpregs_21__30_), .S(n10764), .Z(n10694) );
  MUX2_X2 U15325 ( .A(n10694), .B(n10693), .S(n10878), .Z(n10695) );
  MUX2_X2 U15326 ( .A(decode_regfile_fpregs_18__30_), .B(
        decode_regfile_fpregs_19__30_), .S(n10772), .Z(n10696) );
  MUX2_X2 U15327 ( .A(decode_regfile_fpregs_16__30_), .B(
        decode_regfile_fpregs_17__30_), .S(n10773), .Z(n10697) );
  MUX2_X2 U15328 ( .A(n10697), .B(n10696), .S(n10868), .Z(n10698) );
  MUX2_X2 U15329 ( .A(n10698), .B(n10695), .S(n10921), .Z(n10699) );
  MUX2_X2 U15330 ( .A(n10699), .B(n10692), .S(n10954), .Z(n10700) );
  MUX2_X2 U15331 ( .A(decode_regfile_fpregs_14__30_), .B(
        decode_regfile_fpregs_15__30_), .S(decode_rs2_0_), .Z(n10701) );
  MUX2_X2 U15332 ( .A(decode_regfile_fpregs_12__30_), .B(
        decode_regfile_fpregs_13__30_), .S(n10765), .Z(n10702) );
  MUX2_X2 U15333 ( .A(n10702), .B(n10701), .S(n10871), .Z(n10703) );
  MUX2_X2 U15334 ( .A(decode_regfile_fpregs_10__30_), .B(
        decode_regfile_fpregs_11__30_), .S(n10766), .Z(n10704) );
  MUX2_X2 U15335 ( .A(decode_regfile_fpregs_8__30_), .B(
        decode_regfile_fpregs_9__30_), .S(n10773), .Z(n10705) );
  MUX2_X2 U15336 ( .A(n10705), .B(n10704), .S(n10876), .Z(n10706) );
  MUX2_X2 U15337 ( .A(n10706), .B(n10703), .S(decode_rs2_2_), .Z(n10707) );
  MUX2_X2 U15338 ( .A(decode_regfile_fpregs_6__30_), .B(
        decode_regfile_fpregs_7__30_), .S(n10764), .Z(n10708) );
  MUX2_X2 U15339 ( .A(decode_regfile_fpregs_4__30_), .B(
        decode_regfile_fpregs_5__30_), .S(n10772), .Z(n10709) );
  MUX2_X2 U15340 ( .A(n10709), .B(n10708), .S(n10877), .Z(n10710) );
  MUX2_X2 U15341 ( .A(decode_regfile_fpregs_2__30_), .B(
        decode_regfile_fpregs_3__30_), .S(n10774), .Z(n10711) );
  MUX2_X2 U15342 ( .A(decode_regfile_fpregs_0__30_), .B(
        decode_regfile_fpregs_1__30_), .S(n10775), .Z(n10712) );
  MUX2_X2 U15343 ( .A(n10712), .B(n10711), .S(n10871), .Z(n10713) );
  MUX2_X2 U15344 ( .A(n10713), .B(n10710), .S(decode_rs2_2_), .Z(n10714) );
  MUX2_X2 U15345 ( .A(n10714), .B(n10707), .S(n10954), .Z(n10715) );
  MUX2_X2 U15346 ( .A(n10715), .B(n10700), .S(n10960), .Z(decode_regfile_N29)
         );
  MUX2_X2 U15347 ( .A(decode_regfile_fpregs_30__31_), .B(
        decode_regfile_fpregs_31__31_), .S(n10746), .Z(n10716) );
  MUX2_X2 U15348 ( .A(decode_regfile_fpregs_28__31_), .B(
        decode_regfile_fpregs_29__31_), .S(n10747), .Z(n10717) );
  MUX2_X2 U15349 ( .A(n10717), .B(n10716), .S(n10863), .Z(n10718) );
  MUX2_X2 U15350 ( .A(decode_regfile_fpregs_26__31_), .B(
        decode_regfile_fpregs_27__31_), .S(n10746), .Z(n10719) );
  MUX2_X2 U15351 ( .A(decode_regfile_fpregs_24__31_), .B(
        decode_regfile_fpregs_25__31_), .S(n10765), .Z(n10720) );
  MUX2_X2 U15352 ( .A(n10720), .B(n10719), .S(n10873), .Z(n10721) );
  MUX2_X2 U15353 ( .A(n10721), .B(n10718), .S(decode_rs2_2_), .Z(n10722) );
  MUX2_X2 U15354 ( .A(decode_regfile_fpregs_22__31_), .B(
        decode_regfile_fpregs_23__31_), .S(decode_rs2_0_), .Z(n10723) );
  MUX2_X2 U15355 ( .A(decode_regfile_fpregs_20__31_), .B(
        decode_regfile_fpregs_21__31_), .S(decode_rs2_0_), .Z(n10724) );
  MUX2_X2 U15356 ( .A(n10724), .B(n10723), .S(decode_rs2_1_), .Z(n10725) );
  MUX2_X2 U15357 ( .A(decode_regfile_fpregs_18__31_), .B(
        decode_regfile_fpregs_19__31_), .S(n10766), .Z(n10726) );
  MUX2_X2 U15358 ( .A(decode_regfile_fpregs_16__31_), .B(
        decode_regfile_fpregs_17__31_), .S(n10774), .Z(n10727) );
  MUX2_X2 U15359 ( .A(n10727), .B(n10726), .S(n10872), .Z(n10728) );
  MUX2_X2 U15360 ( .A(n10728), .B(n10725), .S(n10921), .Z(n10729) );
  MUX2_X2 U15361 ( .A(n10729), .B(n10722), .S(n10954), .Z(n10730) );
  MUX2_X2 U15362 ( .A(decode_regfile_fpregs_14__31_), .B(
        decode_regfile_fpregs_15__31_), .S(n10776), .Z(n10731) );
  MUX2_X2 U15363 ( .A(decode_regfile_fpregs_12__31_), .B(
        decode_regfile_fpregs_13__31_), .S(n10764), .Z(n10732) );
  MUX2_X2 U15364 ( .A(n10732), .B(n10731), .S(n10863), .Z(n10733) );
  MUX2_X2 U15365 ( .A(decode_regfile_fpregs_10__31_), .B(
        decode_regfile_fpregs_11__31_), .S(n10772), .Z(n10734) );
  MUX2_X2 U15366 ( .A(decode_regfile_fpregs_8__31_), .B(
        decode_regfile_fpregs_9__31_), .S(n10775), .Z(n10735) );
  MUX2_X2 U15367 ( .A(n10735), .B(n10734), .S(n10878), .Z(n10736) );
  MUX2_X2 U15368 ( .A(n10736), .B(n10733), .S(decode_rs2_2_), .Z(n10737) );
  MUX2_X2 U15369 ( .A(decode_regfile_fpregs_6__31_), .B(
        decode_regfile_fpregs_7__31_), .S(n10765), .Z(n10738) );
  MUX2_X2 U15370 ( .A(decode_regfile_fpregs_4__31_), .B(
        decode_regfile_fpregs_5__31_), .S(n10773), .Z(n10739) );
  MUX2_X2 U15371 ( .A(n10739), .B(n10738), .S(n10875), .Z(n10740) );
  MUX2_X2 U15372 ( .A(decode_regfile_fpregs_2__31_), .B(
        decode_regfile_fpregs_3__31_), .S(n10769), .Z(n10741) );
  MUX2_X2 U15373 ( .A(decode_regfile_fpregs_0__31_), .B(
        decode_regfile_fpregs_1__31_), .S(n10770), .Z(n10742) );
  MUX2_X2 U15374 ( .A(n10742), .B(n10741), .S(n10874), .Z(n10743) );
  MUX2_X2 U15375 ( .A(n10743), .B(n10740), .S(n10921), .Z(n10744) );
  MUX2_X2 U15376 ( .A(n10744), .B(n10737), .S(n10954), .Z(n10745) );
  MUX2_X2 U15377 ( .A(n10745), .B(n10730), .S(n10960), .Z(decode_regfile_N28)
         );
  MUX2_X2 U15378 ( .A(decode_regfile_intregs_28__0_), .B(
        decode_regfile_intregs_29__0_), .S(n12913), .Z(n10962) );
  MUX2_X2 U15379 ( .A(n10962), .B(n10961), .S(n13021), .Z(n10963) );
  MUX2_X2 U15380 ( .A(decode_regfile_intregs_26__0_), .B(
        decode_regfile_intregs_27__0_), .S(n12913), .Z(n10964) );
  MUX2_X2 U15381 ( .A(decode_regfile_intregs_24__0_), .B(
        decode_regfile_intregs_25__0_), .S(n12913), .Z(n10965) );
  MUX2_X2 U15382 ( .A(n10965), .B(n10964), .S(n13021), .Z(n10966) );
  MUX2_X2 U15383 ( .A(n10966), .B(n10963), .S(n13061), .Z(n10967) );
  MUX2_X2 U15384 ( .A(decode_regfile_intregs_22__0_), .B(
        decode_regfile_intregs_23__0_), .S(n12913), .Z(n10968) );
  MUX2_X2 U15385 ( .A(decode_regfile_intregs_20__0_), .B(
        decode_regfile_intregs_21__0_), .S(n12913), .Z(n10969) );
  MUX2_X2 U15386 ( .A(n10969), .B(n10968), .S(n13021), .Z(n10970) );
  MUX2_X2 U15387 ( .A(decode_regfile_intregs_18__0_), .B(
        decode_regfile_intregs_19__0_), .S(n12913), .Z(n10971) );
  MUX2_X2 U15388 ( .A(decode_regfile_intregs_16__0_), .B(
        decode_regfile_intregs_17__0_), .S(n12913), .Z(n10972) );
  MUX2_X2 U15389 ( .A(n10972), .B(n10971), .S(n13021), .Z(n10973) );
  MUX2_X2 U15390 ( .A(n10973), .B(n10970), .S(n13061), .Z(n10974) );
  MUX2_X2 U15391 ( .A(n10974), .B(n10967), .S(decode_rs1_3_), .Z(n10975) );
  MUX2_X2 U15392 ( .A(decode_regfile_intregs_14__0_), .B(
        decode_regfile_intregs_15__0_), .S(n12913), .Z(n10976) );
  MUX2_X2 U15393 ( .A(decode_regfile_intregs_12__0_), .B(
        decode_regfile_intregs_13__0_), .S(n12913), .Z(n10977) );
  MUX2_X2 U15394 ( .A(n10977), .B(n10976), .S(n13021), .Z(n10978) );
  MUX2_X2 U15395 ( .A(decode_regfile_intregs_10__0_), .B(
        decode_regfile_intregs_11__0_), .S(n12913), .Z(n10979) );
  MUX2_X2 U15396 ( .A(decode_regfile_intregs_8__0_), .B(
        decode_regfile_intregs_9__0_), .S(n12913), .Z(n10980) );
  MUX2_X2 U15397 ( .A(n10980), .B(n10979), .S(n13021), .Z(n10981) );
  MUX2_X2 U15398 ( .A(n10981), .B(n10978), .S(n13061), .Z(n10982) );
  MUX2_X2 U15399 ( .A(decode_regfile_intregs_6__0_), .B(
        decode_regfile_intregs_7__0_), .S(n12914), .Z(n10983) );
  MUX2_X2 U15400 ( .A(decode_regfile_intregs_4__0_), .B(
        decode_regfile_intregs_5__0_), .S(n12914), .Z(n10984) );
  MUX2_X2 U15401 ( .A(n10984), .B(n10983), .S(n13022), .Z(n10985) );
  MUX2_X2 U15402 ( .A(decode_regfile_intregs_2__0_), .B(
        decode_regfile_intregs_3__0_), .S(n12914), .Z(n10986) );
  MUX2_X2 U15403 ( .A(decode_regfile_intregs_0__0_), .B(
        decode_regfile_intregs_1__0_), .S(n12914), .Z(n10987) );
  MUX2_X2 U15404 ( .A(n10987), .B(n10986), .S(n13022), .Z(n10988) );
  MUX2_X2 U15405 ( .A(n10988), .B(n10985), .S(n13062), .Z(n10989) );
  MUX2_X2 U15406 ( .A(n10989), .B(n10982), .S(decode_rs1_3_), .Z(n10990) );
  MUX2_X2 U15407 ( .A(n10990), .B(n10975), .S(decode_rs1_4_), .Z(
        decode_regfile_N131) );
  MUX2_X2 U15408 ( .A(decode_regfile_intregs_30__1_), .B(
        decode_regfile_intregs_31__1_), .S(n12914), .Z(n10991) );
  MUX2_X2 U15409 ( .A(decode_regfile_intregs_28__1_), .B(
        decode_regfile_intregs_29__1_), .S(n12914), .Z(n10992) );
  MUX2_X2 U15410 ( .A(n10992), .B(n10991), .S(n13022), .Z(n10993) );
  MUX2_X2 U15411 ( .A(decode_regfile_intregs_26__1_), .B(
        decode_regfile_intregs_27__1_), .S(n12914), .Z(n10994) );
  MUX2_X2 U15412 ( .A(decode_regfile_intregs_24__1_), .B(
        decode_regfile_intregs_25__1_), .S(n12914), .Z(n10995) );
  MUX2_X2 U15413 ( .A(n10995), .B(n10994), .S(n13022), .Z(n10996) );
  MUX2_X2 U15414 ( .A(n10996), .B(n10993), .S(n13062), .Z(n10997) );
  MUX2_X2 U15415 ( .A(decode_regfile_intregs_22__1_), .B(
        decode_regfile_intregs_23__1_), .S(n12914), .Z(n10998) );
  MUX2_X2 U15416 ( .A(decode_regfile_intregs_20__1_), .B(
        decode_regfile_intregs_21__1_), .S(n12914), .Z(n10999) );
  MUX2_X2 U15417 ( .A(n10999), .B(n10998), .S(n13022), .Z(n11000) );
  MUX2_X2 U15418 ( .A(decode_regfile_intregs_18__1_), .B(
        decode_regfile_intregs_19__1_), .S(n12914), .Z(n11001) );
  MUX2_X2 U15419 ( .A(decode_regfile_intregs_16__1_), .B(
        decode_regfile_intregs_17__1_), .S(n12915), .Z(n11002) );
  MUX2_X2 U15420 ( .A(n11002), .B(n11001), .S(n13022), .Z(n11003) );
  MUX2_X2 U15421 ( .A(n11003), .B(n11000), .S(n13062), .Z(n11004) );
  MUX2_X2 U15422 ( .A(n11004), .B(n10997), .S(decode_rs1_3_), .Z(n11005) );
  MUX2_X2 U15423 ( .A(decode_regfile_intregs_14__1_), .B(
        decode_regfile_intregs_15__1_), .S(n12915), .Z(n11006) );
  MUX2_X2 U15424 ( .A(decode_regfile_intregs_12__1_), .B(
        decode_regfile_intregs_13__1_), .S(n12915), .Z(n11007) );
  MUX2_X2 U15425 ( .A(n11007), .B(n11006), .S(n13022), .Z(n11008) );
  MUX2_X2 U15426 ( .A(decode_regfile_intregs_10__1_), .B(
        decode_regfile_intregs_11__1_), .S(n12915), .Z(n11009) );
  MUX2_X2 U15427 ( .A(decode_regfile_intregs_8__1_), .B(
        decode_regfile_intregs_9__1_), .S(n12915), .Z(n11010) );
  MUX2_X2 U15428 ( .A(n11010), .B(n11009), .S(n13022), .Z(n11011) );
  MUX2_X2 U15429 ( .A(n11011), .B(n11008), .S(n13062), .Z(n11012) );
  MUX2_X2 U15430 ( .A(decode_regfile_intregs_6__1_), .B(
        decode_regfile_intregs_7__1_), .S(n12915), .Z(n11013) );
  MUX2_X2 U15431 ( .A(decode_regfile_intregs_4__1_), .B(
        decode_regfile_intregs_5__1_), .S(n12915), .Z(n11014) );
  MUX2_X2 U15432 ( .A(n11014), .B(n11013), .S(n13022), .Z(n11015) );
  MUX2_X2 U15433 ( .A(decode_regfile_intregs_2__1_), .B(
        decode_regfile_intregs_3__1_), .S(n12915), .Z(n11016) );
  MUX2_X2 U15434 ( .A(decode_regfile_intregs_0__1_), .B(
        decode_regfile_intregs_1__1_), .S(n12915), .Z(n11017) );
  MUX2_X2 U15435 ( .A(n11017), .B(n11016), .S(n13022), .Z(n11018) );
  MUX2_X2 U15436 ( .A(n11018), .B(n11015), .S(n13062), .Z(n11019) );
  MUX2_X2 U15437 ( .A(n11019), .B(n11012), .S(decode_rs1_3_), .Z(n11020) );
  MUX2_X2 U15438 ( .A(n11020), .B(n11005), .S(decode_rs1_4_), .Z(
        decode_regfile_N130) );
  MUX2_X2 U15439 ( .A(decode_regfile_intregs_30__2_), .B(
        decode_regfile_intregs_31__2_), .S(n12915), .Z(n11021) );
  MUX2_X2 U15440 ( .A(decode_regfile_intregs_28__2_), .B(
        decode_regfile_intregs_29__2_), .S(n12915), .Z(n11022) );
  MUX2_X2 U15441 ( .A(n11022), .B(n11021), .S(n13022), .Z(n11023) );
  MUX2_X2 U15442 ( .A(decode_regfile_intregs_26__2_), .B(
        decode_regfile_intregs_27__2_), .S(n12916), .Z(n11024) );
  MUX2_X2 U15443 ( .A(decode_regfile_intregs_24__2_), .B(
        decode_regfile_intregs_25__2_), .S(n12916), .Z(n11025) );
  MUX2_X2 U15444 ( .A(n11025), .B(n11024), .S(n13023), .Z(n11026) );
  MUX2_X2 U15445 ( .A(n11026), .B(n11023), .S(n13062), .Z(n11027) );
  MUX2_X2 U15446 ( .A(decode_regfile_intregs_22__2_), .B(
        decode_regfile_intregs_23__2_), .S(n12916), .Z(n11028) );
  MUX2_X2 U15447 ( .A(decode_regfile_intregs_20__2_), .B(
        decode_regfile_intregs_21__2_), .S(n12916), .Z(n11029) );
  MUX2_X2 U15448 ( .A(n11029), .B(n11028), .S(n13023), .Z(n11030) );
  MUX2_X2 U15449 ( .A(decode_regfile_intregs_18__2_), .B(
        decode_regfile_intregs_19__2_), .S(n12916), .Z(n11031) );
  MUX2_X2 U15450 ( .A(decode_regfile_intregs_16__2_), .B(
        decode_regfile_intregs_17__2_), .S(n12916), .Z(n11032) );
  MUX2_X2 U15451 ( .A(n11032), .B(n11031), .S(n13023), .Z(n11033) );
  MUX2_X2 U15452 ( .A(n11033), .B(n11030), .S(n13062), .Z(n11034) );
  MUX2_X2 U15453 ( .A(n11034), .B(n11027), .S(decode_rs1_3_), .Z(n11035) );
  MUX2_X2 U15454 ( .A(decode_regfile_intregs_14__2_), .B(
        decode_regfile_intregs_15__2_), .S(n12916), .Z(n11036) );
  MUX2_X2 U15455 ( .A(decode_regfile_intregs_12__2_), .B(
        decode_regfile_intregs_13__2_), .S(n12916), .Z(n11037) );
  MUX2_X2 U15456 ( .A(n11037), .B(n11036), .S(n13023), .Z(n11038) );
  MUX2_X2 U15457 ( .A(decode_regfile_intregs_10__2_), .B(
        decode_regfile_intregs_11__2_), .S(n12916), .Z(n11039) );
  MUX2_X2 U15458 ( .A(decode_regfile_intregs_8__2_), .B(
        decode_regfile_intregs_9__2_), .S(n12916), .Z(n11040) );
  MUX2_X2 U15459 ( .A(n11040), .B(n11039), .S(n13023), .Z(n11041) );
  MUX2_X2 U15460 ( .A(n11041), .B(n11038), .S(n13062), .Z(n11042) );
  MUX2_X2 U15461 ( .A(decode_regfile_intregs_6__2_), .B(
        decode_regfile_intregs_7__2_), .S(n12916), .Z(n11043) );
  MUX2_X2 U15462 ( .A(decode_regfile_intregs_4__2_), .B(
        decode_regfile_intregs_5__2_), .S(n12917), .Z(n11044) );
  MUX2_X2 U15463 ( .A(n11044), .B(n11043), .S(n13023), .Z(n11045) );
  MUX2_X2 U15464 ( .A(decode_regfile_intregs_2__2_), .B(
        decode_regfile_intregs_3__2_), .S(n12917), .Z(n11046) );
  MUX2_X2 U15465 ( .A(decode_regfile_intregs_0__2_), .B(
        decode_regfile_intregs_1__2_), .S(n12917), .Z(n11047) );
  MUX2_X2 U15466 ( .A(n11047), .B(n11046), .S(n13023), .Z(n11048) );
  MUX2_X2 U15467 ( .A(n11048), .B(n11045), .S(n13062), .Z(n11049) );
  MUX2_X2 U15468 ( .A(n11049), .B(n11042), .S(decode_rs1_3_), .Z(n11050) );
  MUX2_X2 U15469 ( .A(n11050), .B(n11035), .S(decode_rs1_4_), .Z(
        decode_regfile_N129) );
  MUX2_X2 U15470 ( .A(decode_regfile_intregs_30__3_), .B(
        decode_regfile_intregs_31__3_), .S(n12917), .Z(n11051) );
  MUX2_X2 U15471 ( .A(decode_regfile_intregs_28__3_), .B(
        decode_regfile_intregs_29__3_), .S(n12917), .Z(n11052) );
  MUX2_X2 U15472 ( .A(n11052), .B(n11051), .S(n13023), .Z(n11053) );
  MUX2_X2 U15473 ( .A(decode_regfile_intregs_26__3_), .B(
        decode_regfile_intregs_27__3_), .S(n12917), .Z(n11054) );
  MUX2_X2 U15474 ( .A(decode_regfile_intregs_24__3_), .B(
        decode_regfile_intregs_25__3_), .S(n12917), .Z(n11055) );
  MUX2_X2 U15475 ( .A(n11055), .B(n11054), .S(n13023), .Z(n11056) );
  MUX2_X2 U15476 ( .A(n11056), .B(n11053), .S(n13062), .Z(n11057) );
  MUX2_X2 U15477 ( .A(decode_regfile_intregs_22__3_), .B(
        decode_regfile_intregs_23__3_), .S(n12917), .Z(n11058) );
  MUX2_X2 U15478 ( .A(decode_regfile_intregs_20__3_), .B(
        decode_regfile_intregs_21__3_), .S(n12917), .Z(n11059) );
  MUX2_X2 U15479 ( .A(n11059), .B(n11058), .S(n13023), .Z(n11060) );
  MUX2_X2 U15480 ( .A(decode_regfile_intregs_18__3_), .B(
        decode_regfile_intregs_19__3_), .S(n12917), .Z(n11061) );
  MUX2_X2 U15481 ( .A(decode_regfile_intregs_16__3_), .B(
        decode_regfile_intregs_17__3_), .S(n12917), .Z(n11062) );
  MUX2_X2 U15482 ( .A(n11062), .B(n11061), .S(n13023), .Z(n11063) );
  MUX2_X2 U15483 ( .A(n11063), .B(n11060), .S(n13062), .Z(n11064) );
  MUX2_X2 U15484 ( .A(n11064), .B(n11057), .S(decode_rs1_3_), .Z(n11065) );
  MUX2_X2 U15485 ( .A(decode_regfile_intregs_14__3_), .B(
        decode_regfile_intregs_15__3_), .S(n12918), .Z(n11066) );
  MUX2_X2 U15486 ( .A(decode_regfile_intregs_12__3_), .B(
        decode_regfile_intregs_13__3_), .S(n12918), .Z(n11067) );
  MUX2_X2 U15487 ( .A(n11067), .B(n11066), .S(n13024), .Z(n11068) );
  MUX2_X2 U15488 ( .A(decode_regfile_intregs_10__3_), .B(
        decode_regfile_intregs_11__3_), .S(n12918), .Z(n11069) );
  MUX2_X2 U15489 ( .A(decode_regfile_intregs_8__3_), .B(
        decode_regfile_intregs_9__3_), .S(n12918), .Z(n11070) );
  MUX2_X2 U15490 ( .A(n11070), .B(n11069), .S(n13024), .Z(n11071) );
  MUX2_X2 U15491 ( .A(n11071), .B(n11068), .S(n13063), .Z(n11072) );
  MUX2_X2 U15492 ( .A(decode_regfile_intregs_6__3_), .B(
        decode_regfile_intregs_7__3_), .S(n12918), .Z(n11073) );
  MUX2_X2 U15493 ( .A(decode_regfile_intregs_4__3_), .B(
        decode_regfile_intregs_5__3_), .S(n12918), .Z(n11074) );
  MUX2_X2 U15494 ( .A(n11074), .B(n11073), .S(n13024), .Z(n11075) );
  MUX2_X2 U15495 ( .A(decode_regfile_intregs_2__3_), .B(
        decode_regfile_intregs_3__3_), .S(n12918), .Z(n11076) );
  MUX2_X2 U15496 ( .A(decode_regfile_intregs_0__3_), .B(
        decode_regfile_intregs_1__3_), .S(n12918), .Z(n11077) );
  MUX2_X2 U15497 ( .A(n11077), .B(n11076), .S(n13024), .Z(n11078) );
  MUX2_X2 U15498 ( .A(n11078), .B(n11075), .S(n13063), .Z(n11079) );
  MUX2_X2 U15499 ( .A(n11079), .B(n11072), .S(n13084), .Z(n11080) );
  MUX2_X2 U15500 ( .A(n11080), .B(n11065), .S(decode_rs1_4_), .Z(
        decode_regfile_N128) );
  MUX2_X2 U15501 ( .A(decode_regfile_intregs_30__4_), .B(
        decode_regfile_intregs_31__4_), .S(n12918), .Z(n11081) );
  MUX2_X2 U15502 ( .A(decode_regfile_intregs_28__4_), .B(
        decode_regfile_intregs_29__4_), .S(n12918), .Z(n11082) );
  MUX2_X2 U15503 ( .A(n11082), .B(n11081), .S(n13024), .Z(n11083) );
  MUX2_X2 U15504 ( .A(decode_regfile_intregs_26__4_), .B(
        decode_regfile_intregs_27__4_), .S(n12918), .Z(n11084) );
  MUX2_X2 U15505 ( .A(decode_regfile_intregs_24__4_), .B(
        decode_regfile_intregs_25__4_), .S(n12919), .Z(n11085) );
  MUX2_X2 U15506 ( .A(n11085), .B(n11084), .S(n13024), .Z(n11086) );
  MUX2_X2 U15507 ( .A(n11086), .B(n11083), .S(n13063), .Z(n11087) );
  MUX2_X2 U15508 ( .A(decode_regfile_intregs_22__4_), .B(
        decode_regfile_intregs_23__4_), .S(n12919), .Z(n11088) );
  MUX2_X2 U15509 ( .A(decode_regfile_intregs_20__4_), .B(
        decode_regfile_intregs_21__4_), .S(n12919), .Z(n11089) );
  MUX2_X2 U15510 ( .A(n11089), .B(n11088), .S(n13024), .Z(n11090) );
  MUX2_X2 U15511 ( .A(decode_regfile_intregs_18__4_), .B(
        decode_regfile_intregs_19__4_), .S(n12919), .Z(n11091) );
  MUX2_X2 U15512 ( .A(decode_regfile_intregs_16__4_), .B(
        decode_regfile_intregs_17__4_), .S(n12919), .Z(n11092) );
  MUX2_X2 U15513 ( .A(n11092), .B(n11091), .S(n13024), .Z(n11093) );
  MUX2_X2 U15514 ( .A(n11093), .B(n11090), .S(n13063), .Z(n11094) );
  MUX2_X2 U15515 ( .A(n11094), .B(n11087), .S(n13084), .Z(n11095) );
  MUX2_X2 U15516 ( .A(decode_regfile_intregs_14__4_), .B(
        decode_regfile_intregs_15__4_), .S(n12919), .Z(n11096) );
  MUX2_X2 U15517 ( .A(decode_regfile_intregs_12__4_), .B(
        decode_regfile_intregs_13__4_), .S(n12919), .Z(n11097) );
  MUX2_X2 U15518 ( .A(n11097), .B(n11096), .S(n13024), .Z(n11098) );
  MUX2_X2 U15519 ( .A(decode_regfile_intregs_10__4_), .B(
        decode_regfile_intregs_11__4_), .S(n12919), .Z(n11099) );
  MUX2_X2 U15520 ( .A(decode_regfile_intregs_8__4_), .B(
        decode_regfile_intregs_9__4_), .S(n12919), .Z(n11100) );
  MUX2_X2 U15521 ( .A(n11100), .B(n11099), .S(n13024), .Z(n11101) );
  MUX2_X2 U15522 ( .A(n11101), .B(n11098), .S(n13063), .Z(n11102) );
  MUX2_X2 U15523 ( .A(decode_regfile_intregs_6__4_), .B(
        decode_regfile_intregs_7__4_), .S(n12919), .Z(n11103) );
  MUX2_X2 U15524 ( .A(decode_regfile_intregs_4__4_), .B(
        decode_regfile_intregs_5__4_), .S(n12919), .Z(n11104) );
  MUX2_X2 U15525 ( .A(n11104), .B(n11103), .S(n13024), .Z(n11105) );
  MUX2_X2 U15526 ( .A(decode_regfile_intregs_2__4_), .B(
        decode_regfile_intregs_3__4_), .S(n12920), .Z(n11106) );
  MUX2_X2 U15527 ( .A(decode_regfile_intregs_0__4_), .B(
        decode_regfile_intregs_1__4_), .S(n12920), .Z(n11107) );
  MUX2_X2 U15528 ( .A(n11107), .B(n11106), .S(n13025), .Z(n11108) );
  MUX2_X2 U15529 ( .A(n11108), .B(n11105), .S(n13063), .Z(n11109) );
  MUX2_X2 U15530 ( .A(n11109), .B(n11102), .S(n13084), .Z(n11110) );
  MUX2_X2 U15531 ( .A(n11110), .B(n11095), .S(decode_rs1_4_), .Z(
        decode_regfile_N127) );
  MUX2_X2 U15532 ( .A(decode_regfile_intregs_30__5_), .B(
        decode_regfile_intregs_31__5_), .S(n12920), .Z(n11111) );
  MUX2_X2 U15533 ( .A(decode_regfile_intregs_28__5_), .B(
        decode_regfile_intregs_29__5_), .S(n12920), .Z(n11112) );
  MUX2_X2 U15534 ( .A(n11112), .B(n11111), .S(n13025), .Z(n11113) );
  MUX2_X2 U15535 ( .A(decode_regfile_intregs_26__5_), .B(
        decode_regfile_intregs_27__5_), .S(n12920), .Z(n11114) );
  MUX2_X2 U15536 ( .A(decode_regfile_intregs_24__5_), .B(
        decode_regfile_intregs_25__5_), .S(n12920), .Z(n11115) );
  MUX2_X2 U15537 ( .A(n11115), .B(n11114), .S(n13025), .Z(n11116) );
  MUX2_X2 U15538 ( .A(n11116), .B(n11113), .S(n13063), .Z(n11117) );
  MUX2_X2 U15539 ( .A(decode_regfile_intregs_22__5_), .B(
        decode_regfile_intregs_23__5_), .S(n12920), .Z(n11118) );
  MUX2_X2 U15540 ( .A(decode_regfile_intregs_20__5_), .B(
        decode_regfile_intregs_21__5_), .S(n12920), .Z(n11119) );
  MUX2_X2 U15541 ( .A(n11119), .B(n11118), .S(n13025), .Z(n11120) );
  MUX2_X2 U15542 ( .A(decode_regfile_intregs_18__5_), .B(
        decode_regfile_intregs_19__5_), .S(n12920), .Z(n11121) );
  MUX2_X2 U15543 ( .A(decode_regfile_intregs_16__5_), .B(
        decode_regfile_intregs_17__5_), .S(n12920), .Z(n11122) );
  MUX2_X2 U15544 ( .A(n11122), .B(n11121), .S(n13025), .Z(n11123) );
  MUX2_X2 U15545 ( .A(n11123), .B(n11120), .S(n13063), .Z(n11124) );
  MUX2_X2 U15546 ( .A(n11124), .B(n11117), .S(n13084), .Z(n11125) );
  MUX2_X2 U15547 ( .A(decode_regfile_intregs_14__5_), .B(
        decode_regfile_intregs_15__5_), .S(n12920), .Z(n11126) );
  MUX2_X2 U15548 ( .A(decode_regfile_intregs_12__5_), .B(
        decode_regfile_intregs_13__5_), .S(n12921), .Z(n11127) );
  MUX2_X2 U15549 ( .A(n11127), .B(n11126), .S(n13025), .Z(n11128) );
  MUX2_X2 U15550 ( .A(decode_regfile_intregs_10__5_), .B(
        decode_regfile_intregs_11__5_), .S(n12921), .Z(n11129) );
  MUX2_X2 U15551 ( .A(decode_regfile_intregs_8__5_), .B(
        decode_regfile_intregs_9__5_), .S(n12921), .Z(n11130) );
  MUX2_X2 U15552 ( .A(n11130), .B(n11129), .S(n13025), .Z(n11131) );
  MUX2_X2 U15553 ( .A(n11131), .B(n11128), .S(n13063), .Z(n11132) );
  MUX2_X2 U15554 ( .A(decode_regfile_intregs_6__5_), .B(
        decode_regfile_intregs_7__5_), .S(n12921), .Z(n11133) );
  MUX2_X2 U15555 ( .A(decode_regfile_intregs_4__5_), .B(
        decode_regfile_intregs_5__5_), .S(n12921), .Z(n11134) );
  MUX2_X2 U15556 ( .A(n11134), .B(n11133), .S(n13025), .Z(n11135) );
  MUX2_X2 U15557 ( .A(decode_regfile_intregs_2__5_), .B(
        decode_regfile_intregs_3__5_), .S(n12921), .Z(n11136) );
  MUX2_X2 U15558 ( .A(decode_regfile_intregs_0__5_), .B(
        decode_regfile_intregs_1__5_), .S(n12921), .Z(n11137) );
  MUX2_X2 U15559 ( .A(n11137), .B(n11136), .S(n13025), .Z(n11138) );
  MUX2_X2 U15560 ( .A(n11138), .B(n11135), .S(n13063), .Z(n11139) );
  MUX2_X2 U15561 ( .A(n11139), .B(n11132), .S(n13084), .Z(n11140) );
  MUX2_X2 U15562 ( .A(n11140), .B(n11125), .S(decode_rs1_4_), .Z(
        decode_regfile_N126) );
  MUX2_X2 U15563 ( .A(decode_regfile_intregs_30__6_), .B(
        decode_regfile_intregs_31__6_), .S(n12921), .Z(n11141) );
  MUX2_X2 U15564 ( .A(decode_regfile_intregs_28__6_), .B(
        decode_regfile_intregs_29__6_), .S(n12921), .Z(n11142) );
  MUX2_X2 U15565 ( .A(n11142), .B(n11141), .S(n13025), .Z(n11143) );
  MUX2_X2 U15566 ( .A(decode_regfile_intregs_26__6_), .B(
        decode_regfile_intregs_27__6_), .S(n12921), .Z(n11144) );
  MUX2_X2 U15567 ( .A(decode_regfile_intregs_24__6_), .B(
        decode_regfile_intregs_25__6_), .S(n12921), .Z(n11145) );
  MUX2_X2 U15568 ( .A(n11145), .B(n11144), .S(n13025), .Z(n11146) );
  MUX2_X2 U15569 ( .A(n11146), .B(n11143), .S(n13063), .Z(n11147) );
  MUX2_X2 U15570 ( .A(decode_regfile_intregs_22__6_), .B(
        decode_regfile_intregs_23__6_), .S(n12922), .Z(n11148) );
  MUX2_X2 U15571 ( .A(decode_regfile_intregs_20__6_), .B(
        decode_regfile_intregs_21__6_), .S(n12922), .Z(n11149) );
  MUX2_X2 U15572 ( .A(n11149), .B(n11148), .S(n13026), .Z(n11150) );
  MUX2_X2 U15573 ( .A(decode_regfile_intregs_18__6_), .B(
        decode_regfile_intregs_19__6_), .S(n12922), .Z(n11151) );
  MUX2_X2 U15574 ( .A(decode_regfile_intregs_16__6_), .B(
        decode_regfile_intregs_17__6_), .S(n12922), .Z(n11152) );
  MUX2_X2 U15575 ( .A(n11152), .B(n11151), .S(n13026), .Z(n11153) );
  MUX2_X2 U15576 ( .A(n11153), .B(n11150), .S(n13064), .Z(n11154) );
  MUX2_X2 U15577 ( .A(n11154), .B(n11147), .S(n13084), .Z(n11155) );
  MUX2_X2 U15578 ( .A(decode_regfile_intregs_14__6_), .B(
        decode_regfile_intregs_15__6_), .S(n12922), .Z(n11156) );
  MUX2_X2 U15579 ( .A(decode_regfile_intregs_12__6_), .B(
        decode_regfile_intregs_13__6_), .S(n12922), .Z(n11157) );
  MUX2_X2 U15580 ( .A(n11157), .B(n11156), .S(n13026), .Z(n11158) );
  MUX2_X2 U15581 ( .A(decode_regfile_intregs_10__6_), .B(
        decode_regfile_intregs_11__6_), .S(n12922), .Z(n11159) );
  MUX2_X2 U15582 ( .A(decode_regfile_intregs_8__6_), .B(
        decode_regfile_intregs_9__6_), .S(n12922), .Z(n11160) );
  MUX2_X2 U15583 ( .A(n11160), .B(n11159), .S(n13026), .Z(n11161) );
  MUX2_X2 U15584 ( .A(n11161), .B(n11158), .S(n13064), .Z(n11162) );
  MUX2_X2 U15585 ( .A(decode_regfile_intregs_6__6_), .B(
        decode_regfile_intregs_7__6_), .S(n12922), .Z(n11163) );
  MUX2_X2 U15586 ( .A(decode_regfile_intregs_4__6_), .B(
        decode_regfile_intregs_5__6_), .S(n12922), .Z(n11164) );
  MUX2_X2 U15587 ( .A(n11164), .B(n11163), .S(n13026), .Z(n11165) );
  MUX2_X2 U15588 ( .A(decode_regfile_intregs_2__6_), .B(
        decode_regfile_intregs_3__6_), .S(n12922), .Z(n11166) );
  MUX2_X2 U15589 ( .A(decode_regfile_intregs_0__6_), .B(
        decode_regfile_intregs_1__6_), .S(n12923), .Z(n11167) );
  MUX2_X2 U15590 ( .A(n11167), .B(n11166), .S(n13026), .Z(n11168) );
  MUX2_X2 U15591 ( .A(n11168), .B(n11165), .S(n13064), .Z(n11169) );
  MUX2_X2 U15592 ( .A(n11169), .B(n11162), .S(n13084), .Z(n11170) );
  MUX2_X2 U15593 ( .A(n11170), .B(n11155), .S(decode_rs1_4_), .Z(
        decode_regfile_N125) );
  MUX2_X2 U15594 ( .A(decode_regfile_intregs_30__7_), .B(
        decode_regfile_intregs_31__7_), .S(n12923), .Z(n11171) );
  MUX2_X2 U15595 ( .A(decode_regfile_intregs_28__7_), .B(
        decode_regfile_intregs_29__7_), .S(n12923), .Z(n11172) );
  MUX2_X2 U15596 ( .A(n11172), .B(n11171), .S(n13026), .Z(n11173) );
  MUX2_X2 U15597 ( .A(decode_regfile_intregs_26__7_), .B(
        decode_regfile_intregs_27__7_), .S(n12923), .Z(n11174) );
  MUX2_X2 U15598 ( .A(decode_regfile_intregs_24__7_), .B(
        decode_regfile_intregs_25__7_), .S(n12923), .Z(n11175) );
  MUX2_X2 U15599 ( .A(n11175), .B(n11174), .S(n13026), .Z(n11176) );
  MUX2_X2 U15600 ( .A(n11176), .B(n11173), .S(n13064), .Z(n11177) );
  MUX2_X2 U15601 ( .A(decode_regfile_intregs_22__7_), .B(
        decode_regfile_intregs_23__7_), .S(n12923), .Z(n11178) );
  MUX2_X2 U15602 ( .A(decode_regfile_intregs_20__7_), .B(
        decode_regfile_intregs_21__7_), .S(n12923), .Z(n11179) );
  MUX2_X2 U15603 ( .A(n11179), .B(n11178), .S(n13026), .Z(n11180) );
  MUX2_X2 U15604 ( .A(decode_regfile_intregs_18__7_), .B(
        decode_regfile_intregs_19__7_), .S(n12923), .Z(n11181) );
  MUX2_X2 U15605 ( .A(decode_regfile_intregs_16__7_), .B(
        decode_regfile_intregs_17__7_), .S(n12923), .Z(n11182) );
  MUX2_X2 U15606 ( .A(n11182), .B(n11181), .S(n13026), .Z(n11183) );
  MUX2_X2 U15607 ( .A(n11183), .B(n11180), .S(n13064), .Z(n11184) );
  MUX2_X2 U15608 ( .A(n11184), .B(n11177), .S(n13084), .Z(n11185) );
  MUX2_X2 U15609 ( .A(decode_regfile_intregs_14__7_), .B(
        decode_regfile_intregs_15__7_), .S(n12923), .Z(n11186) );
  MUX2_X2 U15610 ( .A(decode_regfile_intregs_12__7_), .B(
        decode_regfile_intregs_13__7_), .S(n12923), .Z(n11187) );
  MUX2_X2 U15611 ( .A(n11187), .B(n11186), .S(n13026), .Z(n11188) );
  MUX2_X2 U15612 ( .A(decode_regfile_intregs_10__7_), .B(
        decode_regfile_intregs_11__7_), .S(n12924), .Z(n11189) );
  MUX2_X2 U15613 ( .A(decode_regfile_intregs_8__7_), .B(
        decode_regfile_intregs_9__7_), .S(n12924), .Z(n11190) );
  MUX2_X2 U15614 ( .A(n11190), .B(n11189), .S(n13027), .Z(n11191) );
  MUX2_X2 U15615 ( .A(n11191), .B(n11188), .S(n13064), .Z(n11192) );
  MUX2_X2 U15616 ( .A(decode_regfile_intregs_6__7_), .B(
        decode_regfile_intregs_7__7_), .S(n12924), .Z(n11193) );
  MUX2_X2 U15617 ( .A(decode_regfile_intregs_4__7_), .B(
        decode_regfile_intregs_5__7_), .S(n12924), .Z(n11194) );
  MUX2_X2 U15618 ( .A(n11194), .B(n11193), .S(n13027), .Z(n11195) );
  MUX2_X2 U15619 ( .A(decode_regfile_intregs_2__7_), .B(
        decode_regfile_intregs_3__7_), .S(n12924), .Z(n11196) );
  MUX2_X2 U15620 ( .A(decode_regfile_intregs_0__7_), .B(
        decode_regfile_intregs_1__7_), .S(n12924), .Z(n11197) );
  MUX2_X2 U15621 ( .A(n11197), .B(n11196), .S(n13027), .Z(n11198) );
  MUX2_X2 U15622 ( .A(n11198), .B(n11195), .S(n13064), .Z(n11199) );
  MUX2_X2 U15623 ( .A(n11199), .B(n11192), .S(n13084), .Z(n11200) );
  MUX2_X2 U15624 ( .A(n11200), .B(n11185), .S(decode_rs1_4_), .Z(
        decode_regfile_N124) );
  MUX2_X2 U15625 ( .A(decode_regfile_intregs_30__8_), .B(
        decode_regfile_intregs_31__8_), .S(n12924), .Z(n11201) );
  MUX2_X2 U15626 ( .A(decode_regfile_intregs_28__8_), .B(
        decode_regfile_intregs_29__8_), .S(n12924), .Z(n11202) );
  MUX2_X2 U15627 ( .A(n11202), .B(n11201), .S(n13027), .Z(n11203) );
  MUX2_X2 U15628 ( .A(decode_regfile_intregs_26__8_), .B(
        decode_regfile_intregs_27__8_), .S(n12924), .Z(n11204) );
  MUX2_X2 U15629 ( .A(decode_regfile_intregs_24__8_), .B(
        decode_regfile_intregs_25__8_), .S(n12924), .Z(n11205) );
  MUX2_X2 U15630 ( .A(n11205), .B(n11204), .S(n13027), .Z(n11206) );
  MUX2_X2 U15631 ( .A(n11206), .B(n11203), .S(n13064), .Z(n11207) );
  MUX2_X2 U15632 ( .A(decode_regfile_intregs_22__8_), .B(
        decode_regfile_intregs_23__8_), .S(n12924), .Z(n11208) );
  MUX2_X2 U15633 ( .A(decode_regfile_intregs_20__8_), .B(
        decode_regfile_intregs_21__8_), .S(n12925), .Z(n11209) );
  MUX2_X2 U15634 ( .A(n11209), .B(n11208), .S(n13027), .Z(n11210) );
  MUX2_X2 U15635 ( .A(decode_regfile_intregs_18__8_), .B(
        decode_regfile_intregs_19__8_), .S(n12925), .Z(n11211) );
  MUX2_X2 U15636 ( .A(decode_regfile_intregs_16__8_), .B(
        decode_regfile_intregs_17__8_), .S(n12925), .Z(n11212) );
  MUX2_X2 U15637 ( .A(n11212), .B(n11211), .S(n13027), .Z(n11213) );
  MUX2_X2 U15638 ( .A(n11213), .B(n11210), .S(n13064), .Z(n11214) );
  MUX2_X2 U15639 ( .A(n11214), .B(n11207), .S(n13084), .Z(n11215) );
  MUX2_X2 U15640 ( .A(decode_regfile_intregs_14__8_), .B(
        decode_regfile_intregs_15__8_), .S(n12925), .Z(n11216) );
  MUX2_X2 U15641 ( .A(decode_regfile_intregs_12__8_), .B(
        decode_regfile_intregs_13__8_), .S(n12925), .Z(n11217) );
  MUX2_X2 U15642 ( .A(n11217), .B(n11216), .S(n13027), .Z(n11218) );
  MUX2_X2 U15643 ( .A(decode_regfile_intregs_10__8_), .B(
        decode_regfile_intregs_11__8_), .S(n12925), .Z(n11219) );
  MUX2_X2 U15644 ( .A(decode_regfile_intregs_8__8_), .B(
        decode_regfile_intregs_9__8_), .S(n12925), .Z(n11220) );
  MUX2_X2 U15645 ( .A(n11220), .B(n11219), .S(n13027), .Z(n11221) );
  MUX2_X2 U15646 ( .A(n11221), .B(n11218), .S(n13064), .Z(n11222) );
  MUX2_X2 U15647 ( .A(decode_regfile_intregs_6__8_), .B(
        decode_regfile_intregs_7__8_), .S(n12925), .Z(n11223) );
  MUX2_X2 U15648 ( .A(decode_regfile_intregs_4__8_), .B(
        decode_regfile_intregs_5__8_), .S(n12925), .Z(n11224) );
  MUX2_X2 U15649 ( .A(n11224), .B(n11223), .S(n13027), .Z(n11225) );
  MUX2_X2 U15650 ( .A(decode_regfile_intregs_2__8_), .B(
        decode_regfile_intregs_3__8_), .S(n12925), .Z(n11226) );
  MUX2_X2 U15651 ( .A(decode_regfile_intregs_0__8_), .B(
        decode_regfile_intregs_1__8_), .S(n12925), .Z(n11227) );
  MUX2_X2 U15652 ( .A(n11227), .B(n11226), .S(n13027), .Z(n11228) );
  MUX2_X2 U15653 ( .A(n11228), .B(n11225), .S(n13064), .Z(n11229) );
  MUX2_X2 U15654 ( .A(n11229), .B(n11222), .S(n13084), .Z(n11230) );
  MUX2_X2 U15655 ( .A(n11230), .B(n11215), .S(decode_rs1_4_), .Z(
        decode_regfile_N123) );
  MUX2_X2 U15656 ( .A(decode_regfile_intregs_30__9_), .B(
        decode_regfile_intregs_31__9_), .S(n12926), .Z(n11231) );
  MUX2_X2 U15657 ( .A(decode_regfile_intregs_28__9_), .B(
        decode_regfile_intregs_29__9_), .S(n12926), .Z(n11232) );
  MUX2_X2 U15658 ( .A(n11232), .B(n11231), .S(n13028), .Z(n11233) );
  MUX2_X2 U15659 ( .A(decode_regfile_intregs_26__9_), .B(
        decode_regfile_intregs_27__9_), .S(n12926), .Z(n11234) );
  MUX2_X2 U15660 ( .A(decode_regfile_intregs_24__9_), .B(
        decode_regfile_intregs_25__9_), .S(n12926), .Z(n11235) );
  MUX2_X2 U15661 ( .A(n11235), .B(n11234), .S(n13028), .Z(n11236) );
  MUX2_X2 U15662 ( .A(n11236), .B(n11233), .S(n13065), .Z(n11237) );
  MUX2_X2 U15663 ( .A(decode_regfile_intregs_22__9_), .B(
        decode_regfile_intregs_23__9_), .S(n12926), .Z(n11238) );
  MUX2_X2 U15664 ( .A(decode_regfile_intregs_20__9_), .B(
        decode_regfile_intregs_21__9_), .S(n12926), .Z(n11239) );
  MUX2_X2 U15665 ( .A(n11239), .B(n11238), .S(n13028), .Z(n11240) );
  MUX2_X2 U15666 ( .A(decode_regfile_intregs_18__9_), .B(
        decode_regfile_intregs_19__9_), .S(n12926), .Z(n11241) );
  MUX2_X2 U15667 ( .A(decode_regfile_intregs_16__9_), .B(
        decode_regfile_intregs_17__9_), .S(n12926), .Z(n11242) );
  MUX2_X2 U15668 ( .A(n11242), .B(n11241), .S(n13028), .Z(n11243) );
  MUX2_X2 U15669 ( .A(n11243), .B(n11240), .S(n13065), .Z(n11244) );
  MUX2_X2 U15670 ( .A(n11244), .B(n11237), .S(n13085), .Z(n11245) );
  MUX2_X2 U15671 ( .A(decode_regfile_intregs_14__9_), .B(
        decode_regfile_intregs_15__9_), .S(n12926), .Z(n11246) );
  MUX2_X2 U15672 ( .A(decode_regfile_intregs_12__9_), .B(
        decode_regfile_intregs_13__9_), .S(n12926), .Z(n11247) );
  MUX2_X2 U15673 ( .A(n11247), .B(n11246), .S(n13028), .Z(n11248) );
  MUX2_X2 U15674 ( .A(decode_regfile_intregs_10__9_), .B(
        decode_regfile_intregs_11__9_), .S(n12926), .Z(n11249) );
  MUX2_X2 U15675 ( .A(decode_regfile_intregs_8__9_), .B(
        decode_regfile_intregs_9__9_), .S(n12927), .Z(n11250) );
  MUX2_X2 U15676 ( .A(n11250), .B(n11249), .S(n13028), .Z(n11251) );
  MUX2_X2 U15677 ( .A(n11251), .B(n11248), .S(n13065), .Z(n11252) );
  MUX2_X2 U15678 ( .A(decode_regfile_intregs_6__9_), .B(
        decode_regfile_intregs_7__9_), .S(n12927), .Z(n11253) );
  MUX2_X2 U15679 ( .A(decode_regfile_intregs_4__9_), .B(
        decode_regfile_intregs_5__9_), .S(n12927), .Z(n11254) );
  MUX2_X2 U15680 ( .A(n11254), .B(n11253), .S(n13028), .Z(n11255) );
  MUX2_X2 U15681 ( .A(decode_regfile_intregs_2__9_), .B(
        decode_regfile_intregs_3__9_), .S(n12927), .Z(n11256) );
  MUX2_X2 U15682 ( .A(decode_regfile_intregs_0__9_), .B(
        decode_regfile_intregs_1__9_), .S(n12927), .Z(n11257) );
  MUX2_X2 U15683 ( .A(n11257), .B(n11256), .S(n13028), .Z(n11258) );
  MUX2_X2 U15684 ( .A(n11258), .B(n11255), .S(n13065), .Z(n11259) );
  MUX2_X2 U15685 ( .A(n11259), .B(n11252), .S(n13085), .Z(n11260) );
  MUX2_X2 U15686 ( .A(n11260), .B(n11245), .S(n13097), .Z(decode_regfile_N122)
         );
  MUX2_X2 U15687 ( .A(decode_regfile_intregs_30__10_), .B(
        decode_regfile_intregs_31__10_), .S(n12927), .Z(n11261) );
  MUX2_X2 U15688 ( .A(decode_regfile_intregs_28__10_), .B(
        decode_regfile_intregs_29__10_), .S(n12927), .Z(n11262) );
  MUX2_X2 U15689 ( .A(n11262), .B(n11261), .S(n13028), .Z(n11263) );
  MUX2_X2 U15690 ( .A(decode_regfile_intregs_26__10_), .B(
        decode_regfile_intregs_27__10_), .S(n12927), .Z(n11264) );
  MUX2_X2 U15691 ( .A(decode_regfile_intregs_24__10_), .B(
        decode_regfile_intregs_25__10_), .S(n12927), .Z(n11265) );
  MUX2_X2 U15692 ( .A(n11265), .B(n11264), .S(n13028), .Z(n11266) );
  MUX2_X2 U15693 ( .A(n11266), .B(n11263), .S(n13065), .Z(n11267) );
  MUX2_X2 U15694 ( .A(decode_regfile_intregs_22__10_), .B(
        decode_regfile_intregs_23__10_), .S(n12927), .Z(n11268) );
  MUX2_X2 U15695 ( .A(decode_regfile_intregs_20__10_), .B(
        decode_regfile_intregs_21__10_), .S(n12927), .Z(n11269) );
  MUX2_X2 U15696 ( .A(n11269), .B(n11268), .S(n13028), .Z(n11270) );
  MUX2_X2 U15697 ( .A(decode_regfile_intregs_18__10_), .B(
        decode_regfile_intregs_19__10_), .S(n12928), .Z(n11271) );
  MUX2_X2 U15698 ( .A(decode_regfile_intregs_16__10_), .B(
        decode_regfile_intregs_17__10_), .S(n12928), .Z(n11272) );
  MUX2_X2 U15699 ( .A(n11272), .B(n11271), .S(n13029), .Z(n11273) );
  MUX2_X2 U15700 ( .A(n11273), .B(n11270), .S(n13065), .Z(n11274) );
  MUX2_X2 U15701 ( .A(n11274), .B(n11267), .S(n13085), .Z(n11275) );
  MUX2_X2 U15702 ( .A(decode_regfile_intregs_14__10_), .B(
        decode_regfile_intregs_15__10_), .S(n12928), .Z(n11276) );
  MUX2_X2 U15703 ( .A(decode_regfile_intregs_12__10_), .B(
        decode_regfile_intregs_13__10_), .S(n12928), .Z(n11277) );
  MUX2_X2 U15704 ( .A(n11277), .B(n11276), .S(n13029), .Z(n11278) );
  MUX2_X2 U15705 ( .A(decode_regfile_intregs_10__10_), .B(
        decode_regfile_intregs_11__10_), .S(n12928), .Z(n11279) );
  MUX2_X2 U15706 ( .A(decode_regfile_intregs_8__10_), .B(
        decode_regfile_intregs_9__10_), .S(n12928), .Z(n11280) );
  MUX2_X2 U15707 ( .A(n11280), .B(n11279), .S(n13029), .Z(n11281) );
  MUX2_X2 U15708 ( .A(n11281), .B(n11278), .S(n13065), .Z(n11282) );
  MUX2_X2 U15709 ( .A(decode_regfile_intregs_6__10_), .B(
        decode_regfile_intregs_7__10_), .S(n12928), .Z(n11283) );
  MUX2_X2 U15710 ( .A(decode_regfile_intregs_4__10_), .B(
        decode_regfile_intregs_5__10_), .S(n12928), .Z(n11284) );
  MUX2_X2 U15711 ( .A(n11284), .B(n11283), .S(n13029), .Z(n11285) );
  MUX2_X2 U15712 ( .A(decode_regfile_intregs_2__10_), .B(
        decode_regfile_intregs_3__10_), .S(n12928), .Z(n11286) );
  MUX2_X2 U15713 ( .A(decode_regfile_intregs_0__10_), .B(
        decode_regfile_intregs_1__10_), .S(n12928), .Z(n11287) );
  MUX2_X2 U15714 ( .A(n11287), .B(n11286), .S(n13029), .Z(n11288) );
  MUX2_X2 U15715 ( .A(n11288), .B(n11285), .S(n13065), .Z(n11289) );
  MUX2_X2 U15716 ( .A(n11289), .B(n11282), .S(n13085), .Z(n11290) );
  MUX2_X2 U15717 ( .A(n11290), .B(n11275), .S(n13097), .Z(decode_regfile_N121)
         );
  MUX2_X2 U15718 ( .A(decode_regfile_intregs_30__11_), .B(
        decode_regfile_intregs_31__11_), .S(n12928), .Z(n11291) );
  MUX2_X2 U15719 ( .A(decode_regfile_intregs_28__11_), .B(
        decode_regfile_intregs_29__11_), .S(n12929), .Z(n11292) );
  MUX2_X2 U15720 ( .A(n11292), .B(n11291), .S(n13029), .Z(n11293) );
  MUX2_X2 U15721 ( .A(decode_regfile_intregs_26__11_), .B(
        decode_regfile_intregs_27__11_), .S(n12929), .Z(n11294) );
  MUX2_X2 U15722 ( .A(decode_regfile_intregs_24__11_), .B(
        decode_regfile_intregs_25__11_), .S(n12929), .Z(n11295) );
  MUX2_X2 U15723 ( .A(n11295), .B(n11294), .S(n13029), .Z(n11296) );
  MUX2_X2 U15724 ( .A(n11296), .B(n11293), .S(n13065), .Z(n11297) );
  MUX2_X2 U15725 ( .A(decode_regfile_intregs_22__11_), .B(
        decode_regfile_intregs_23__11_), .S(n12929), .Z(n11298) );
  MUX2_X2 U15726 ( .A(decode_regfile_intregs_20__11_), .B(
        decode_regfile_intregs_21__11_), .S(n12929), .Z(n11299) );
  MUX2_X2 U15727 ( .A(n11299), .B(n11298), .S(n13029), .Z(n11300) );
  MUX2_X2 U15728 ( .A(decode_regfile_intregs_18__11_), .B(
        decode_regfile_intregs_19__11_), .S(n12929), .Z(n11301) );
  MUX2_X2 U15729 ( .A(decode_regfile_intregs_16__11_), .B(
        decode_regfile_intregs_17__11_), .S(n12929), .Z(n11302) );
  MUX2_X2 U15730 ( .A(n11302), .B(n11301), .S(n13029), .Z(n11303) );
  MUX2_X2 U15731 ( .A(n11303), .B(n11300), .S(n13065), .Z(n11304) );
  MUX2_X2 U15732 ( .A(n11304), .B(n11297), .S(n13085), .Z(n11305) );
  MUX2_X2 U15733 ( .A(decode_regfile_intregs_14__11_), .B(
        decode_regfile_intregs_15__11_), .S(n12929), .Z(n11306) );
  MUX2_X2 U15734 ( .A(decode_regfile_intregs_12__11_), .B(
        decode_regfile_intregs_13__11_), .S(n12929), .Z(n11307) );
  MUX2_X2 U15735 ( .A(n11307), .B(n11306), .S(n13029), .Z(n11308) );
  MUX2_X2 U15736 ( .A(decode_regfile_intregs_10__11_), .B(
        decode_regfile_intregs_11__11_), .S(n12929), .Z(n11309) );
  MUX2_X2 U15737 ( .A(decode_regfile_intregs_8__11_), .B(
        decode_regfile_intregs_9__11_), .S(n12929), .Z(n11310) );
  MUX2_X2 U15738 ( .A(n11310), .B(n11309), .S(n13029), .Z(n11311) );
  MUX2_X2 U15739 ( .A(n11311), .B(n11308), .S(n13065), .Z(n11312) );
  MUX2_X2 U15740 ( .A(decode_regfile_intregs_6__11_), .B(
        decode_regfile_intregs_7__11_), .S(n12930), .Z(n11313) );
  MUX2_X2 U15741 ( .A(decode_regfile_intregs_4__11_), .B(
        decode_regfile_intregs_5__11_), .S(n12930), .Z(n11314) );
  MUX2_X2 U15742 ( .A(n11314), .B(n11313), .S(n13030), .Z(n11315) );
  MUX2_X2 U15743 ( .A(decode_regfile_intregs_2__11_), .B(
        decode_regfile_intregs_3__11_), .S(n12930), .Z(n11316) );
  MUX2_X2 U15744 ( .A(decode_regfile_intregs_0__11_), .B(
        decode_regfile_intregs_1__11_), .S(n12930), .Z(n11317) );
  MUX2_X2 U15745 ( .A(n11317), .B(n11316), .S(n13030), .Z(n11318) );
  MUX2_X2 U15746 ( .A(n11318), .B(n11315), .S(n13066), .Z(n11319) );
  MUX2_X2 U15747 ( .A(n11319), .B(n11312), .S(n13085), .Z(n11320) );
  MUX2_X2 U15748 ( .A(n11320), .B(n11305), .S(n13097), .Z(decode_regfile_N120)
         );
  MUX2_X2 U15749 ( .A(decode_regfile_intregs_30__12_), .B(
        decode_regfile_intregs_31__12_), .S(n12930), .Z(n11321) );
  MUX2_X2 U15750 ( .A(decode_regfile_intregs_28__12_), .B(
        decode_regfile_intregs_29__12_), .S(n12930), .Z(n11322) );
  MUX2_X2 U15751 ( .A(n11322), .B(n11321), .S(n13030), .Z(n11323) );
  MUX2_X2 U15752 ( .A(decode_regfile_intregs_26__12_), .B(
        decode_regfile_intregs_27__12_), .S(n12930), .Z(n11324) );
  MUX2_X2 U15753 ( .A(decode_regfile_intregs_24__12_), .B(
        decode_regfile_intregs_25__12_), .S(n12930), .Z(n11325) );
  MUX2_X2 U15754 ( .A(n11325), .B(n11324), .S(n13030), .Z(n11326) );
  MUX2_X2 U15755 ( .A(n11326), .B(n11323), .S(n13066), .Z(n11327) );
  MUX2_X2 U15756 ( .A(decode_regfile_intregs_22__12_), .B(
        decode_regfile_intregs_23__12_), .S(n12930), .Z(n11328) );
  MUX2_X2 U15757 ( .A(decode_regfile_intregs_20__12_), .B(
        decode_regfile_intregs_21__12_), .S(n12930), .Z(n11329) );
  MUX2_X2 U15758 ( .A(n11329), .B(n11328), .S(n13030), .Z(n11330) );
  MUX2_X2 U15759 ( .A(decode_regfile_intregs_18__12_), .B(
        decode_regfile_intregs_19__12_), .S(n12930), .Z(n11331) );
  MUX2_X2 U15760 ( .A(decode_regfile_intregs_16__12_), .B(
        decode_regfile_intregs_17__12_), .S(n12931), .Z(n11332) );
  MUX2_X2 U15761 ( .A(n11332), .B(n11331), .S(n13030), .Z(n11333) );
  MUX2_X2 U15762 ( .A(n11333), .B(n11330), .S(n13066), .Z(n11334) );
  MUX2_X2 U15763 ( .A(n11334), .B(n11327), .S(n13085), .Z(n11335) );
  MUX2_X2 U15764 ( .A(decode_regfile_intregs_14__12_), .B(
        decode_regfile_intregs_15__12_), .S(n12931), .Z(n11336) );
  MUX2_X2 U15765 ( .A(decode_regfile_intregs_12__12_), .B(
        decode_regfile_intregs_13__12_), .S(n12931), .Z(n11337) );
  MUX2_X2 U15766 ( .A(n11337), .B(n11336), .S(n13030), .Z(n11338) );
  MUX2_X2 U15767 ( .A(decode_regfile_intregs_10__12_), .B(
        decode_regfile_intregs_11__12_), .S(n12931), .Z(n11339) );
  MUX2_X2 U15768 ( .A(decode_regfile_intregs_8__12_), .B(
        decode_regfile_intregs_9__12_), .S(n12931), .Z(n11340) );
  MUX2_X2 U15769 ( .A(n11340), .B(n11339), .S(n13030), .Z(n11341) );
  MUX2_X2 U15770 ( .A(n11341), .B(n11338), .S(n13066), .Z(n11342) );
  MUX2_X2 U15771 ( .A(decode_regfile_intregs_6__12_), .B(
        decode_regfile_intregs_7__12_), .S(n12931), .Z(n11343) );
  MUX2_X2 U15772 ( .A(decode_regfile_intregs_4__12_), .B(
        decode_regfile_intregs_5__12_), .S(n12931), .Z(n11344) );
  MUX2_X2 U15773 ( .A(n11344), .B(n11343), .S(n13030), .Z(n11345) );
  MUX2_X2 U15774 ( .A(decode_regfile_intregs_2__12_), .B(
        decode_regfile_intregs_3__12_), .S(n12931), .Z(n11346) );
  MUX2_X2 U15775 ( .A(decode_regfile_intregs_0__12_), .B(
        decode_regfile_intregs_1__12_), .S(n12931), .Z(n11347) );
  MUX2_X2 U15776 ( .A(n11347), .B(n11346), .S(n13030), .Z(n11348) );
  MUX2_X2 U15777 ( .A(n11348), .B(n11345), .S(n13066), .Z(n11349) );
  MUX2_X2 U15778 ( .A(n11349), .B(n11342), .S(n13085), .Z(n11350) );
  MUX2_X2 U15779 ( .A(n11350), .B(n11335), .S(n13097), .Z(decode_regfile_N119)
         );
  MUX2_X2 U15780 ( .A(decode_regfile_intregs_30__13_), .B(
        decode_regfile_intregs_31__13_), .S(n12931), .Z(n11351) );
  MUX2_X2 U15781 ( .A(decode_regfile_intregs_28__13_), .B(
        decode_regfile_intregs_29__13_), .S(n12931), .Z(n11352) );
  MUX2_X2 U15782 ( .A(n11352), .B(n11351), .S(n13030), .Z(n11353) );
  MUX2_X2 U15783 ( .A(decode_regfile_intregs_26__13_), .B(
        decode_regfile_intregs_27__13_), .S(n12932), .Z(n11354) );
  MUX2_X2 U15784 ( .A(decode_regfile_intregs_24__13_), .B(
        decode_regfile_intregs_25__13_), .S(n12932), .Z(n11355) );
  MUX2_X2 U15785 ( .A(n11355), .B(n11354), .S(n13031), .Z(n11356) );
  MUX2_X2 U15786 ( .A(n11356), .B(n11353), .S(n13066), .Z(n11357) );
  MUX2_X2 U15787 ( .A(decode_regfile_intregs_22__13_), .B(
        decode_regfile_intregs_23__13_), .S(n12932), .Z(n11358) );
  MUX2_X2 U15788 ( .A(decode_regfile_intregs_20__13_), .B(
        decode_regfile_intregs_21__13_), .S(n12932), .Z(n11359) );
  MUX2_X2 U15789 ( .A(n11359), .B(n11358), .S(n13031), .Z(n11360) );
  MUX2_X2 U15790 ( .A(decode_regfile_intregs_18__13_), .B(
        decode_regfile_intregs_19__13_), .S(n12932), .Z(n11361) );
  MUX2_X2 U15791 ( .A(decode_regfile_intregs_16__13_), .B(
        decode_regfile_intregs_17__13_), .S(n12932), .Z(n11362) );
  MUX2_X2 U15792 ( .A(n11362), .B(n11361), .S(n13031), .Z(n11363) );
  MUX2_X2 U15793 ( .A(n11363), .B(n11360), .S(n13066), .Z(n11364) );
  MUX2_X2 U15794 ( .A(n11364), .B(n11357), .S(n13085), .Z(n11365) );
  MUX2_X2 U15795 ( .A(decode_regfile_intregs_14__13_), .B(
        decode_regfile_intregs_15__13_), .S(n12932), .Z(n11366) );
  MUX2_X2 U15796 ( .A(decode_regfile_intregs_12__13_), .B(
        decode_regfile_intregs_13__13_), .S(n12932), .Z(n11367) );
  MUX2_X2 U15797 ( .A(n11367), .B(n11366), .S(n13031), .Z(n11368) );
  MUX2_X2 U15798 ( .A(decode_regfile_intregs_10__13_), .B(
        decode_regfile_intregs_11__13_), .S(n12932), .Z(n11369) );
  MUX2_X2 U15799 ( .A(decode_regfile_intregs_8__13_), .B(
        decode_regfile_intregs_9__13_), .S(n12932), .Z(n11370) );
  MUX2_X2 U15800 ( .A(n11370), .B(n11369), .S(n13031), .Z(n11371) );
  MUX2_X2 U15801 ( .A(n11371), .B(n11368), .S(n13066), .Z(n11372) );
  MUX2_X2 U15802 ( .A(decode_regfile_intregs_6__13_), .B(
        decode_regfile_intregs_7__13_), .S(n12932), .Z(n11373) );
  MUX2_X2 U15803 ( .A(decode_regfile_intregs_4__13_), .B(
        decode_regfile_intregs_5__13_), .S(n12933), .Z(n11374) );
  MUX2_X2 U15804 ( .A(n11374), .B(n11373), .S(n13031), .Z(n11375) );
  MUX2_X2 U15805 ( .A(decode_regfile_intregs_2__13_), .B(
        decode_regfile_intregs_3__13_), .S(n12933), .Z(n11376) );
  MUX2_X2 U15806 ( .A(decode_regfile_intregs_0__13_), .B(
        decode_regfile_intregs_1__13_), .S(n12933), .Z(n11377) );
  MUX2_X2 U15807 ( .A(n11377), .B(n11376), .S(n13031), .Z(n11378) );
  MUX2_X2 U15808 ( .A(n11378), .B(n11375), .S(n13066), .Z(n11379) );
  MUX2_X2 U15809 ( .A(n11379), .B(n11372), .S(n13085), .Z(n11380) );
  MUX2_X2 U15810 ( .A(n11380), .B(n11365), .S(n13097), .Z(decode_regfile_N118)
         );
  MUX2_X2 U15811 ( .A(decode_regfile_intregs_30__14_), .B(
        decode_regfile_intregs_31__14_), .S(n12933), .Z(n11381) );
  MUX2_X2 U15812 ( .A(decode_regfile_intregs_28__14_), .B(
        decode_regfile_intregs_29__14_), .S(n12933), .Z(n11382) );
  MUX2_X2 U15813 ( .A(n11382), .B(n11381), .S(n13031), .Z(n11383) );
  MUX2_X2 U15814 ( .A(decode_regfile_intregs_26__14_), .B(
        decode_regfile_intregs_27__14_), .S(n12933), .Z(n11384) );
  MUX2_X2 U15815 ( .A(decode_regfile_intregs_24__14_), .B(
        decode_regfile_intregs_25__14_), .S(n12933), .Z(n11385) );
  MUX2_X2 U15816 ( .A(n11385), .B(n11384), .S(n13031), .Z(n11386) );
  MUX2_X2 U15817 ( .A(n11386), .B(n11383), .S(n13066), .Z(n11387) );
  MUX2_X2 U15818 ( .A(decode_regfile_intregs_22__14_), .B(
        decode_regfile_intregs_23__14_), .S(n12933), .Z(n11388) );
  MUX2_X2 U15819 ( .A(decode_regfile_intregs_20__14_), .B(
        decode_regfile_intregs_21__14_), .S(n12933), .Z(n11389) );
  MUX2_X2 U15820 ( .A(n11389), .B(n11388), .S(n13031), .Z(n11390) );
  MUX2_X2 U15821 ( .A(decode_regfile_intregs_18__14_), .B(
        decode_regfile_intregs_19__14_), .S(n12933), .Z(n11391) );
  MUX2_X2 U15822 ( .A(decode_regfile_intregs_16__14_), .B(
        decode_regfile_intregs_17__14_), .S(n12933), .Z(n11392) );
  MUX2_X2 U15823 ( .A(n11392), .B(n11391), .S(n13031), .Z(n11393) );
  MUX2_X2 U15824 ( .A(n11393), .B(n11390), .S(n13066), .Z(n11394) );
  MUX2_X2 U15825 ( .A(n11394), .B(n11387), .S(n13085), .Z(n11395) );
  MUX2_X2 U15826 ( .A(decode_regfile_intregs_14__14_), .B(
        decode_regfile_intregs_15__14_), .S(n12934), .Z(n11396) );
  MUX2_X2 U15827 ( .A(decode_regfile_intregs_12__14_), .B(
        decode_regfile_intregs_13__14_), .S(n12934), .Z(n11397) );
  MUX2_X2 U15828 ( .A(n11397), .B(n11396), .S(n13032), .Z(n11398) );
  MUX2_X2 U15829 ( .A(decode_regfile_intregs_10__14_), .B(
        decode_regfile_intregs_11__14_), .S(n12934), .Z(n11399) );
  MUX2_X2 U15830 ( .A(decode_regfile_intregs_8__14_), .B(
        decode_regfile_intregs_9__14_), .S(n12934), .Z(n11400) );
  MUX2_X2 U15831 ( .A(n11400), .B(n11399), .S(n13032), .Z(n11401) );
  MUX2_X2 U15832 ( .A(n11401), .B(n11398), .S(n13067), .Z(n11402) );
  MUX2_X2 U15833 ( .A(decode_regfile_intregs_6__14_), .B(
        decode_regfile_intregs_7__14_), .S(n12934), .Z(n11403) );
  MUX2_X2 U15834 ( .A(decode_regfile_intregs_4__14_), .B(
        decode_regfile_intregs_5__14_), .S(n12934), .Z(n11404) );
  MUX2_X2 U15835 ( .A(n11404), .B(n11403), .S(n13032), .Z(n11405) );
  MUX2_X2 U15836 ( .A(decode_regfile_intregs_2__14_), .B(
        decode_regfile_intregs_3__14_), .S(n12934), .Z(n11406) );
  MUX2_X2 U15837 ( .A(decode_regfile_intregs_0__14_), .B(
        decode_regfile_intregs_1__14_), .S(n12934), .Z(n11407) );
  MUX2_X2 U15838 ( .A(n11407), .B(n11406), .S(n13032), .Z(n11408) );
  MUX2_X2 U15839 ( .A(n11408), .B(n11405), .S(n13067), .Z(n11409) );
  MUX2_X2 U15840 ( .A(n11409), .B(n11402), .S(n13086), .Z(n11410) );
  MUX2_X2 U15841 ( .A(n11410), .B(n11395), .S(n13097), .Z(decode_regfile_N117)
         );
  MUX2_X2 U15842 ( .A(decode_regfile_intregs_30__15_), .B(
        decode_regfile_intregs_31__15_), .S(n12934), .Z(n11411) );
  MUX2_X2 U15843 ( .A(decode_regfile_intregs_28__15_), .B(
        decode_regfile_intregs_29__15_), .S(n12934), .Z(n11412) );
  MUX2_X2 U15844 ( .A(n11412), .B(n11411), .S(n13032), .Z(n11413) );
  MUX2_X2 U15845 ( .A(decode_regfile_intregs_26__15_), .B(
        decode_regfile_intregs_27__15_), .S(n12934), .Z(n11414) );
  MUX2_X2 U15846 ( .A(decode_regfile_intregs_24__15_), .B(
        decode_regfile_intregs_25__15_), .S(n12935), .Z(n11415) );
  MUX2_X2 U15847 ( .A(n11415), .B(n11414), .S(n13032), .Z(n11416) );
  MUX2_X2 U15848 ( .A(n11416), .B(n11413), .S(n13067), .Z(n11417) );
  MUX2_X2 U15849 ( .A(decode_regfile_intregs_22__15_), .B(
        decode_regfile_intregs_23__15_), .S(n12935), .Z(n11418) );
  MUX2_X2 U15850 ( .A(decode_regfile_intregs_20__15_), .B(
        decode_regfile_intregs_21__15_), .S(n12935), .Z(n11419) );
  MUX2_X2 U15851 ( .A(n11419), .B(n11418), .S(n13032), .Z(n11420) );
  MUX2_X2 U15852 ( .A(decode_regfile_intregs_18__15_), .B(
        decode_regfile_intregs_19__15_), .S(n12935), .Z(n11421) );
  MUX2_X2 U15853 ( .A(decode_regfile_intregs_16__15_), .B(
        decode_regfile_intregs_17__15_), .S(n12935), .Z(n11422) );
  MUX2_X2 U15854 ( .A(n11422), .B(n11421), .S(n13032), .Z(n11423) );
  MUX2_X2 U15855 ( .A(n11423), .B(n11420), .S(n13067), .Z(n11424) );
  MUX2_X2 U15856 ( .A(n11424), .B(n11417), .S(n13086), .Z(n11425) );
  MUX2_X2 U15857 ( .A(decode_regfile_intregs_14__15_), .B(
        decode_regfile_intregs_15__15_), .S(n12935), .Z(n11426) );
  MUX2_X2 U15858 ( .A(decode_regfile_intregs_12__15_), .B(
        decode_regfile_intregs_13__15_), .S(n12935), .Z(n11427) );
  MUX2_X2 U15859 ( .A(n11427), .B(n11426), .S(n13032), .Z(n11428) );
  MUX2_X2 U15860 ( .A(decode_regfile_intregs_10__15_), .B(
        decode_regfile_intregs_11__15_), .S(n12935), .Z(n11429) );
  MUX2_X2 U15861 ( .A(decode_regfile_intregs_8__15_), .B(
        decode_regfile_intregs_9__15_), .S(n12935), .Z(n11430) );
  MUX2_X2 U15862 ( .A(n11430), .B(n11429), .S(n13032), .Z(n11431) );
  MUX2_X2 U15863 ( .A(n11431), .B(n11428), .S(n13067), .Z(n11432) );
  MUX2_X2 U15864 ( .A(decode_regfile_intregs_6__15_), .B(
        decode_regfile_intregs_7__15_), .S(n12935), .Z(n11433) );
  MUX2_X2 U15865 ( .A(decode_regfile_intregs_4__15_), .B(
        decode_regfile_intregs_5__15_), .S(n12935), .Z(n11434) );
  MUX2_X2 U15866 ( .A(n11434), .B(n11433), .S(n13032), .Z(n11435) );
  MUX2_X2 U15867 ( .A(decode_regfile_intregs_2__15_), .B(
        decode_regfile_intregs_3__15_), .S(n12936), .Z(n11436) );
  MUX2_X2 U15868 ( .A(decode_regfile_intregs_0__15_), .B(
        decode_regfile_intregs_1__15_), .S(n12936), .Z(n11437) );
  MUX2_X2 U15869 ( .A(n11437), .B(n11436), .S(n13033), .Z(n11438) );
  MUX2_X2 U15870 ( .A(n11438), .B(n11435), .S(n13067), .Z(n11439) );
  MUX2_X2 U15871 ( .A(n11439), .B(n11432), .S(n13086), .Z(n11440) );
  MUX2_X2 U15872 ( .A(n11440), .B(n11425), .S(n13097), .Z(decode_regfile_N116)
         );
  MUX2_X2 U15873 ( .A(decode_regfile_intregs_30__16_), .B(
        decode_regfile_intregs_31__16_), .S(n12936), .Z(n11441) );
  MUX2_X2 U15874 ( .A(decode_regfile_intregs_28__16_), .B(
        decode_regfile_intregs_29__16_), .S(n12936), .Z(n11442) );
  MUX2_X2 U15875 ( .A(n11442), .B(n11441), .S(n13033), .Z(n11443) );
  MUX2_X2 U15876 ( .A(decode_regfile_intregs_26__16_), .B(
        decode_regfile_intregs_27__16_), .S(n12936), .Z(n11444) );
  MUX2_X2 U15877 ( .A(decode_regfile_intregs_24__16_), .B(
        decode_regfile_intregs_25__16_), .S(n12936), .Z(n11445) );
  MUX2_X2 U15878 ( .A(n11445), .B(n11444), .S(n13033), .Z(n11446) );
  MUX2_X2 U15879 ( .A(n11446), .B(n11443), .S(n13067), .Z(n11447) );
  MUX2_X2 U15880 ( .A(decode_regfile_intregs_22__16_), .B(
        decode_regfile_intregs_23__16_), .S(n12936), .Z(n11448) );
  MUX2_X2 U15881 ( .A(decode_regfile_intregs_20__16_), .B(
        decode_regfile_intregs_21__16_), .S(n12936), .Z(n11449) );
  MUX2_X2 U15882 ( .A(n11449), .B(n11448), .S(n13033), .Z(n11450) );
  MUX2_X2 U15883 ( .A(decode_regfile_intregs_18__16_), .B(
        decode_regfile_intregs_19__16_), .S(n12936), .Z(n11451) );
  MUX2_X2 U15884 ( .A(decode_regfile_intregs_16__16_), .B(
        decode_regfile_intregs_17__16_), .S(n12936), .Z(n11452) );
  MUX2_X2 U15885 ( .A(n11452), .B(n11451), .S(n13033), .Z(n11453) );
  MUX2_X2 U15886 ( .A(n11453), .B(n11450), .S(n13067), .Z(n11454) );
  MUX2_X2 U15887 ( .A(n11454), .B(n11447), .S(n13086), .Z(n11455) );
  MUX2_X2 U15888 ( .A(decode_regfile_intregs_14__16_), .B(
        decode_regfile_intregs_15__16_), .S(n12936), .Z(n11456) );
  MUX2_X2 U15889 ( .A(decode_regfile_intregs_12__16_), .B(
        decode_regfile_intregs_13__16_), .S(n12937), .Z(n11457) );
  MUX2_X2 U15890 ( .A(n11457), .B(n11456), .S(n13033), .Z(n11458) );
  MUX2_X2 U15891 ( .A(decode_regfile_intregs_10__16_), .B(
        decode_regfile_intregs_11__16_), .S(n12937), .Z(n11459) );
  MUX2_X2 U15892 ( .A(decode_regfile_intregs_8__16_), .B(
        decode_regfile_intregs_9__16_), .S(n12937), .Z(n11460) );
  MUX2_X2 U15893 ( .A(n11460), .B(n11459), .S(n13033), .Z(n11461) );
  MUX2_X2 U15894 ( .A(n11461), .B(n11458), .S(n13067), .Z(n11462) );
  MUX2_X2 U15895 ( .A(decode_regfile_intregs_6__16_), .B(
        decode_regfile_intregs_7__16_), .S(n12937), .Z(n11463) );
  MUX2_X2 U15896 ( .A(decode_regfile_intregs_4__16_), .B(
        decode_regfile_intregs_5__16_), .S(n12937), .Z(n11464) );
  MUX2_X2 U15897 ( .A(n11464), .B(n11463), .S(n13033), .Z(n11465) );
  MUX2_X2 U15898 ( .A(decode_regfile_intregs_2__16_), .B(
        decode_regfile_intregs_3__16_), .S(n12937), .Z(n11466) );
  MUX2_X2 U15899 ( .A(decode_regfile_intregs_0__16_), .B(
        decode_regfile_intregs_1__16_), .S(n12937), .Z(n11467) );
  MUX2_X2 U15900 ( .A(n11467), .B(n11466), .S(n13033), .Z(n11468) );
  MUX2_X2 U15901 ( .A(n11468), .B(n11465), .S(n13067), .Z(n11469) );
  MUX2_X2 U15902 ( .A(n11469), .B(n11462), .S(n13086), .Z(n11470) );
  MUX2_X2 U15903 ( .A(n11470), .B(n11455), .S(n13097), .Z(decode_regfile_N115)
         );
  MUX2_X2 U15904 ( .A(decode_regfile_intregs_30__17_), .B(
        decode_regfile_intregs_31__17_), .S(n12937), .Z(n11471) );
  MUX2_X2 U15905 ( .A(decode_regfile_intregs_28__17_), .B(
        decode_regfile_intregs_29__17_), .S(n12937), .Z(n11472) );
  MUX2_X2 U15906 ( .A(n11472), .B(n11471), .S(n13033), .Z(n11473) );
  MUX2_X2 U15907 ( .A(decode_regfile_intregs_26__17_), .B(
        decode_regfile_intregs_27__17_), .S(n12937), .Z(n11474) );
  MUX2_X2 U15908 ( .A(decode_regfile_intregs_24__17_), .B(
        decode_regfile_intregs_25__17_), .S(n12937), .Z(n11475) );
  MUX2_X2 U15909 ( .A(n11475), .B(n11474), .S(n13033), .Z(n11476) );
  MUX2_X2 U15910 ( .A(n11476), .B(n11473), .S(n13067), .Z(n11477) );
  MUX2_X2 U15911 ( .A(decode_regfile_intregs_22__17_), .B(
        decode_regfile_intregs_23__17_), .S(n12938), .Z(n11478) );
  MUX2_X2 U15912 ( .A(decode_regfile_intregs_20__17_), .B(
        decode_regfile_intregs_21__17_), .S(n12938), .Z(n11479) );
  MUX2_X2 U15913 ( .A(n11479), .B(n11478), .S(n13034), .Z(n11480) );
  MUX2_X2 U15914 ( .A(decode_regfile_intregs_18__17_), .B(
        decode_regfile_intregs_19__17_), .S(n12938), .Z(n11481) );
  MUX2_X2 U15915 ( .A(decode_regfile_intregs_16__17_), .B(
        decode_regfile_intregs_17__17_), .S(n12938), .Z(n11482) );
  MUX2_X2 U15916 ( .A(n11482), .B(n11481), .S(n13034), .Z(n11483) );
  MUX2_X2 U15917 ( .A(n11483), .B(n11480), .S(n13068), .Z(n11484) );
  MUX2_X2 U15918 ( .A(n11484), .B(n11477), .S(n13086), .Z(n11485) );
  MUX2_X2 U15919 ( .A(decode_regfile_intregs_14__17_), .B(
        decode_regfile_intregs_15__17_), .S(n12938), .Z(n11486) );
  MUX2_X2 U15920 ( .A(decode_regfile_intregs_12__17_), .B(
        decode_regfile_intregs_13__17_), .S(n12938), .Z(n11487) );
  MUX2_X2 U15921 ( .A(n11487), .B(n11486), .S(n13034), .Z(n11488) );
  MUX2_X2 U15922 ( .A(decode_regfile_intregs_10__17_), .B(
        decode_regfile_intregs_11__17_), .S(n12938), .Z(n11489) );
  MUX2_X2 U15923 ( .A(decode_regfile_intregs_8__17_), .B(
        decode_regfile_intregs_9__17_), .S(n12938), .Z(n11490) );
  MUX2_X2 U15924 ( .A(n11490), .B(n11489), .S(n13034), .Z(n11491) );
  MUX2_X2 U15925 ( .A(n11491), .B(n11488), .S(n13068), .Z(n11492) );
  MUX2_X2 U15926 ( .A(decode_regfile_intregs_6__17_), .B(
        decode_regfile_intregs_7__17_), .S(n12938), .Z(n11493) );
  MUX2_X2 U15927 ( .A(decode_regfile_intregs_4__17_), .B(
        decode_regfile_intregs_5__17_), .S(n12938), .Z(n11494) );
  MUX2_X2 U15928 ( .A(n11494), .B(n11493), .S(n13034), .Z(n11495) );
  MUX2_X2 U15929 ( .A(decode_regfile_intregs_2__17_), .B(
        decode_regfile_intregs_3__17_), .S(n12938), .Z(n11496) );
  MUX2_X2 U15930 ( .A(decode_regfile_intregs_0__17_), .B(
        decode_regfile_intregs_1__17_), .S(n12939), .Z(n11497) );
  MUX2_X2 U15931 ( .A(n11497), .B(n11496), .S(n13034), .Z(n11498) );
  MUX2_X2 U15932 ( .A(n11498), .B(n11495), .S(n13068), .Z(n11499) );
  MUX2_X2 U15933 ( .A(n11499), .B(n11492), .S(n13086), .Z(n11500) );
  MUX2_X2 U15934 ( .A(n11500), .B(n11485), .S(n13097), .Z(decode_regfile_N114)
         );
  MUX2_X2 U15935 ( .A(decode_regfile_intregs_30__18_), .B(
        decode_regfile_intregs_31__18_), .S(n12939), .Z(n11501) );
  MUX2_X2 U15936 ( .A(decode_regfile_intregs_28__18_), .B(
        decode_regfile_intregs_29__18_), .S(n12939), .Z(n11502) );
  MUX2_X2 U15937 ( .A(n11502), .B(n11501), .S(n13034), .Z(n11503) );
  MUX2_X2 U15938 ( .A(decode_regfile_intregs_26__18_), .B(
        decode_regfile_intregs_27__18_), .S(n12939), .Z(n11504) );
  MUX2_X2 U15939 ( .A(decode_regfile_intregs_24__18_), .B(
        decode_regfile_intregs_25__18_), .S(n12939), .Z(n11505) );
  MUX2_X2 U15940 ( .A(n11505), .B(n11504), .S(n13034), .Z(n11506) );
  MUX2_X2 U15941 ( .A(n11506), .B(n11503), .S(n13068), .Z(n11507) );
  MUX2_X2 U15942 ( .A(decode_regfile_intregs_22__18_), .B(
        decode_regfile_intregs_23__18_), .S(n12939), .Z(n11508) );
  MUX2_X2 U15943 ( .A(decode_regfile_intregs_20__18_), .B(
        decode_regfile_intregs_21__18_), .S(n12939), .Z(n11509) );
  MUX2_X2 U15944 ( .A(n11509), .B(n11508), .S(n13034), .Z(n11510) );
  MUX2_X2 U15945 ( .A(decode_regfile_intregs_18__18_), .B(
        decode_regfile_intregs_19__18_), .S(n12939), .Z(n11511) );
  MUX2_X2 U15946 ( .A(decode_regfile_intregs_16__18_), .B(
        decode_regfile_intregs_17__18_), .S(n12939), .Z(n11512) );
  MUX2_X2 U15947 ( .A(n11512), .B(n11511), .S(n13034), .Z(n11513) );
  MUX2_X2 U15948 ( .A(n11513), .B(n11510), .S(n13068), .Z(n11514) );
  MUX2_X2 U15949 ( .A(n11514), .B(n11507), .S(n13086), .Z(n11515) );
  MUX2_X2 U15950 ( .A(decode_regfile_intregs_14__18_), .B(
        decode_regfile_intregs_15__18_), .S(n12939), .Z(n11516) );
  MUX2_X2 U15951 ( .A(decode_regfile_intregs_12__18_), .B(
        decode_regfile_intregs_13__18_), .S(n12939), .Z(n11517) );
  MUX2_X2 U15952 ( .A(n11517), .B(n11516), .S(n13034), .Z(n11518) );
  MUX2_X2 U15953 ( .A(decode_regfile_intregs_10__18_), .B(
        decode_regfile_intregs_11__18_), .S(n12940), .Z(n11519) );
  MUX2_X2 U15954 ( .A(decode_regfile_intregs_8__18_), .B(
        decode_regfile_intregs_9__18_), .S(n12940), .Z(n11520) );
  MUX2_X2 U15955 ( .A(n11520), .B(n11519), .S(n13035), .Z(n11521) );
  MUX2_X2 U15956 ( .A(n11521), .B(n11518), .S(n13068), .Z(n11522) );
  MUX2_X2 U15957 ( .A(decode_regfile_intregs_6__18_), .B(
        decode_regfile_intregs_7__18_), .S(n12940), .Z(n11523) );
  MUX2_X2 U15958 ( .A(decode_regfile_intregs_4__18_), .B(
        decode_regfile_intregs_5__18_), .S(n12940), .Z(n11524) );
  MUX2_X2 U15959 ( .A(n11524), .B(n11523), .S(n13035), .Z(n11525) );
  MUX2_X2 U15960 ( .A(decode_regfile_intregs_2__18_), .B(
        decode_regfile_intregs_3__18_), .S(n12940), .Z(n11526) );
  MUX2_X2 U15961 ( .A(decode_regfile_intregs_0__18_), .B(
        decode_regfile_intregs_1__18_), .S(n12940), .Z(n11527) );
  MUX2_X2 U15962 ( .A(n11527), .B(n11526), .S(n13035), .Z(n11528) );
  MUX2_X2 U15963 ( .A(n11528), .B(n11525), .S(n13068), .Z(n11529) );
  MUX2_X2 U15964 ( .A(n11529), .B(n11522), .S(n13086), .Z(n11530) );
  MUX2_X2 U15965 ( .A(n11530), .B(n11515), .S(n13097), .Z(decode_regfile_N113)
         );
  MUX2_X2 U15966 ( .A(decode_regfile_intregs_30__19_), .B(
        decode_regfile_intregs_31__19_), .S(n12940), .Z(n11531) );
  MUX2_X2 U15967 ( .A(decode_regfile_intregs_28__19_), .B(
        decode_regfile_intregs_29__19_), .S(n12940), .Z(n11532) );
  MUX2_X2 U15968 ( .A(n11532), .B(n11531), .S(n13035), .Z(n11533) );
  MUX2_X2 U15969 ( .A(decode_regfile_intregs_26__19_), .B(
        decode_regfile_intregs_27__19_), .S(n12940), .Z(n11534) );
  MUX2_X2 U15970 ( .A(decode_regfile_intregs_24__19_), .B(
        decode_regfile_intregs_25__19_), .S(n12940), .Z(n11535) );
  MUX2_X2 U15971 ( .A(n11535), .B(n11534), .S(n13035), .Z(n11536) );
  MUX2_X2 U15972 ( .A(n11536), .B(n11533), .S(n13068), .Z(n11537) );
  MUX2_X2 U15973 ( .A(decode_regfile_intregs_22__19_), .B(
        decode_regfile_intregs_23__19_), .S(n12940), .Z(n11538) );
  MUX2_X2 U15974 ( .A(decode_regfile_intregs_20__19_), .B(
        decode_regfile_intregs_21__19_), .S(n12941), .Z(n11539) );
  MUX2_X2 U15975 ( .A(n11539), .B(n11538), .S(n13035), .Z(n11540) );
  MUX2_X2 U15976 ( .A(decode_regfile_intregs_18__19_), .B(
        decode_regfile_intregs_19__19_), .S(n12941), .Z(n11541) );
  MUX2_X2 U15977 ( .A(decode_regfile_intregs_16__19_), .B(
        decode_regfile_intregs_17__19_), .S(n12941), .Z(n11542) );
  MUX2_X2 U15978 ( .A(n11542), .B(n11541), .S(n13035), .Z(n11543) );
  MUX2_X2 U15979 ( .A(n11543), .B(n11540), .S(n13068), .Z(n11544) );
  MUX2_X2 U15980 ( .A(n11544), .B(n11537), .S(n13086), .Z(n11545) );
  MUX2_X2 U15981 ( .A(decode_regfile_intregs_14__19_), .B(
        decode_regfile_intregs_15__19_), .S(n12941), .Z(n11546) );
  MUX2_X2 U15982 ( .A(decode_regfile_intregs_12__19_), .B(
        decode_regfile_intregs_13__19_), .S(n12941), .Z(n11547) );
  MUX2_X2 U15983 ( .A(n11547), .B(n11546), .S(n13035), .Z(n11548) );
  MUX2_X2 U15984 ( .A(decode_regfile_intregs_10__19_), .B(
        decode_regfile_intregs_11__19_), .S(n12941), .Z(n11549) );
  MUX2_X2 U15985 ( .A(decode_regfile_intregs_8__19_), .B(
        decode_regfile_intregs_9__19_), .S(n12941), .Z(n11550) );
  MUX2_X2 U15986 ( .A(n11550), .B(n11549), .S(n13035), .Z(n11551) );
  MUX2_X2 U15987 ( .A(n11551), .B(n11548), .S(n13068), .Z(n11552) );
  MUX2_X2 U15988 ( .A(decode_regfile_intregs_6__19_), .B(
        decode_regfile_intregs_7__19_), .S(n12941), .Z(n11553) );
  MUX2_X2 U15989 ( .A(decode_regfile_intregs_4__19_), .B(
        decode_regfile_intregs_5__19_), .S(n12941), .Z(n11554) );
  MUX2_X2 U15990 ( .A(n11554), .B(n11553), .S(n13035), .Z(n11555) );
  MUX2_X2 U15991 ( .A(decode_regfile_intregs_2__19_), .B(
        decode_regfile_intregs_3__19_), .S(n12941), .Z(n11556) );
  MUX2_X2 U15992 ( .A(decode_regfile_intregs_0__19_), .B(
        decode_regfile_intregs_1__19_), .S(n12941), .Z(n11557) );
  MUX2_X2 U15993 ( .A(n11557), .B(n11556), .S(n13035), .Z(n11558) );
  MUX2_X2 U15994 ( .A(n11558), .B(n11555), .S(n13068), .Z(n11559) );
  MUX2_X2 U15995 ( .A(n11559), .B(n11552), .S(n13086), .Z(n11560) );
  MUX2_X2 U15996 ( .A(n11560), .B(n11545), .S(n13097), .Z(decode_regfile_N112)
         );
  MUX2_X2 U15997 ( .A(decode_regfile_intregs_30__20_), .B(
        decode_regfile_intregs_31__20_), .S(n12942), .Z(n11561) );
  MUX2_X2 U15998 ( .A(decode_regfile_intregs_28__20_), .B(
        decode_regfile_intregs_29__20_), .S(n12942), .Z(n11562) );
  MUX2_X2 U15999 ( .A(n11562), .B(n11561), .S(n13036), .Z(n11563) );
  MUX2_X2 U16000 ( .A(decode_regfile_intregs_26__20_), .B(
        decode_regfile_intregs_27__20_), .S(n12942), .Z(n11564) );
  MUX2_X2 U16001 ( .A(decode_regfile_intregs_24__20_), .B(
        decode_regfile_intregs_25__20_), .S(n12942), .Z(n11565) );
  MUX2_X2 U16002 ( .A(n11565), .B(n11564), .S(n13036), .Z(n11566) );
  MUX2_X2 U16003 ( .A(n11566), .B(n11563), .S(n13069), .Z(n11567) );
  MUX2_X2 U16004 ( .A(decode_regfile_intregs_22__20_), .B(
        decode_regfile_intregs_23__20_), .S(n12942), .Z(n11568) );
  MUX2_X2 U16005 ( .A(decode_regfile_intregs_20__20_), .B(
        decode_regfile_intregs_21__20_), .S(n12942), .Z(n11569) );
  MUX2_X2 U16006 ( .A(n11569), .B(n11568), .S(n13036), .Z(n11570) );
  MUX2_X2 U16007 ( .A(decode_regfile_intregs_18__20_), .B(
        decode_regfile_intregs_19__20_), .S(n12942), .Z(n11571) );
  MUX2_X2 U16008 ( .A(decode_regfile_intregs_16__20_), .B(
        decode_regfile_intregs_17__20_), .S(n12942), .Z(n11572) );
  MUX2_X2 U16009 ( .A(n11572), .B(n11571), .S(n13036), .Z(n11573) );
  MUX2_X2 U16010 ( .A(n11573), .B(n11570), .S(n13069), .Z(n11574) );
  MUX2_X2 U16011 ( .A(n11574), .B(n11567), .S(n13087), .Z(n11575) );
  MUX2_X2 U16012 ( .A(decode_regfile_intregs_14__20_), .B(
        decode_regfile_intregs_15__20_), .S(n12942), .Z(n11576) );
  MUX2_X2 U16013 ( .A(decode_regfile_intregs_12__20_), .B(
        decode_regfile_intregs_13__20_), .S(n12942), .Z(n11577) );
  MUX2_X2 U16014 ( .A(n11577), .B(n11576), .S(n13036), .Z(n11578) );
  MUX2_X2 U16015 ( .A(decode_regfile_intregs_10__20_), .B(
        decode_regfile_intregs_11__20_), .S(n12942), .Z(n11579) );
  MUX2_X2 U16016 ( .A(decode_regfile_intregs_8__20_), .B(
        decode_regfile_intregs_9__20_), .S(n12943), .Z(n11580) );
  MUX2_X2 U16017 ( .A(n11580), .B(n11579), .S(n13036), .Z(n11581) );
  MUX2_X2 U16018 ( .A(n11581), .B(n11578), .S(n13069), .Z(n11582) );
  MUX2_X2 U16019 ( .A(decode_regfile_intregs_6__20_), .B(
        decode_regfile_intregs_7__20_), .S(n12943), .Z(n11583) );
  MUX2_X2 U16020 ( .A(decode_regfile_intregs_4__20_), .B(
        decode_regfile_intregs_5__20_), .S(n12943), .Z(n11584) );
  MUX2_X2 U16021 ( .A(n11584), .B(n11583), .S(n13036), .Z(n11585) );
  MUX2_X2 U16022 ( .A(decode_regfile_intregs_2__20_), .B(
        decode_regfile_intregs_3__20_), .S(n12943), .Z(n11586) );
  MUX2_X2 U16023 ( .A(decode_regfile_intregs_0__20_), .B(
        decode_regfile_intregs_1__20_), .S(n12943), .Z(n11587) );
  MUX2_X2 U16024 ( .A(n11587), .B(n11586), .S(n13036), .Z(n11588) );
  MUX2_X2 U16025 ( .A(n11588), .B(n11585), .S(n13069), .Z(n11589) );
  MUX2_X2 U16026 ( .A(n11589), .B(n11582), .S(n13087), .Z(n11590) );
  MUX2_X2 U16027 ( .A(n11590), .B(n11575), .S(n13098), .Z(decode_regfile_N111)
         );
  MUX2_X2 U16028 ( .A(decode_regfile_intregs_30__21_), .B(
        decode_regfile_intregs_31__21_), .S(n12943), .Z(n11591) );
  MUX2_X2 U16029 ( .A(decode_regfile_intregs_28__21_), .B(
        decode_regfile_intregs_29__21_), .S(n12943), .Z(n11592) );
  MUX2_X2 U16030 ( .A(n11592), .B(n11591), .S(n13036), .Z(n11593) );
  MUX2_X2 U16031 ( .A(decode_regfile_intregs_26__21_), .B(
        decode_regfile_intregs_27__21_), .S(n12943), .Z(n11594) );
  MUX2_X2 U16032 ( .A(decode_regfile_intregs_24__21_), .B(
        decode_regfile_intregs_25__21_), .S(n12943), .Z(n11595) );
  MUX2_X2 U16033 ( .A(n11595), .B(n11594), .S(n13036), .Z(n11596) );
  MUX2_X2 U16034 ( .A(n11596), .B(n11593), .S(n13069), .Z(n11597) );
  MUX2_X2 U16035 ( .A(decode_regfile_intregs_22__21_), .B(
        decode_regfile_intregs_23__21_), .S(n12943), .Z(n11598) );
  MUX2_X2 U16036 ( .A(decode_regfile_intregs_20__21_), .B(
        decode_regfile_intregs_21__21_), .S(n12943), .Z(n11599) );
  MUX2_X2 U16037 ( .A(n11599), .B(n11598), .S(n13036), .Z(n11600) );
  MUX2_X2 U16038 ( .A(decode_regfile_intregs_18__21_), .B(
        decode_regfile_intregs_19__21_), .S(n12944), .Z(n11601) );
  MUX2_X2 U16039 ( .A(decode_regfile_intregs_16__21_), .B(
        decode_regfile_intregs_17__21_), .S(n12944), .Z(n11602) );
  MUX2_X2 U16040 ( .A(n11602), .B(n11601), .S(n13037), .Z(n11603) );
  MUX2_X2 U16041 ( .A(n11603), .B(n11600), .S(n13069), .Z(n11604) );
  MUX2_X2 U16042 ( .A(n11604), .B(n11597), .S(n13087), .Z(n11605) );
  MUX2_X2 U16043 ( .A(decode_regfile_intregs_14__21_), .B(
        decode_regfile_intregs_15__21_), .S(n12944), .Z(n11606) );
  MUX2_X2 U16044 ( .A(decode_regfile_intregs_12__21_), .B(
        decode_regfile_intregs_13__21_), .S(n12944), .Z(n11607) );
  MUX2_X2 U16045 ( .A(n11607), .B(n11606), .S(n13037), .Z(n11608) );
  MUX2_X2 U16046 ( .A(decode_regfile_intregs_10__21_), .B(
        decode_regfile_intregs_11__21_), .S(n12944), .Z(n11609) );
  MUX2_X2 U16047 ( .A(decode_regfile_intregs_8__21_), .B(
        decode_regfile_intregs_9__21_), .S(n12944), .Z(n11610) );
  MUX2_X2 U16048 ( .A(n11610), .B(n11609), .S(n13037), .Z(n11611) );
  MUX2_X2 U16049 ( .A(n11611), .B(n11608), .S(n13069), .Z(n11612) );
  MUX2_X2 U16050 ( .A(decode_regfile_intregs_6__21_), .B(
        decode_regfile_intregs_7__21_), .S(n12944), .Z(n11613) );
  MUX2_X2 U16051 ( .A(decode_regfile_intregs_4__21_), .B(
        decode_regfile_intregs_5__21_), .S(n12944), .Z(n11614) );
  MUX2_X2 U16052 ( .A(n11614), .B(n11613), .S(n13037), .Z(n11615) );
  MUX2_X2 U16053 ( .A(decode_regfile_intregs_2__21_), .B(
        decode_regfile_intregs_3__21_), .S(n12944), .Z(n11616) );
  MUX2_X2 U16054 ( .A(decode_regfile_intregs_0__21_), .B(
        decode_regfile_intregs_1__21_), .S(n12944), .Z(n11617) );
  MUX2_X2 U16055 ( .A(n11617), .B(n11616), .S(n13037), .Z(n11618) );
  MUX2_X2 U16056 ( .A(n11618), .B(n11615), .S(n13069), .Z(n11619) );
  MUX2_X2 U16057 ( .A(n11619), .B(n11612), .S(n13087), .Z(n11620) );
  MUX2_X2 U16058 ( .A(n11620), .B(n11605), .S(n13098), .Z(decode_regfile_N110)
         );
  MUX2_X2 U16059 ( .A(decode_regfile_intregs_30__22_), .B(
        decode_regfile_intregs_31__22_), .S(n12944), .Z(n11621) );
  MUX2_X2 U16060 ( .A(decode_regfile_intregs_28__22_), .B(
        decode_regfile_intregs_29__22_), .S(n12945), .Z(n11622) );
  MUX2_X2 U16061 ( .A(n11622), .B(n11621), .S(n13037), .Z(n11623) );
  MUX2_X2 U16062 ( .A(decode_regfile_intregs_26__22_), .B(
        decode_regfile_intregs_27__22_), .S(n12945), .Z(n11624) );
  MUX2_X2 U16063 ( .A(decode_regfile_intregs_24__22_), .B(
        decode_regfile_intregs_25__22_), .S(n12945), .Z(n11625) );
  MUX2_X2 U16064 ( .A(n11625), .B(n11624), .S(n13037), .Z(n11626) );
  MUX2_X2 U16065 ( .A(n11626), .B(n11623), .S(n13069), .Z(n11627) );
  MUX2_X2 U16066 ( .A(decode_regfile_intregs_22__22_), .B(
        decode_regfile_intregs_23__22_), .S(n12945), .Z(n11628) );
  MUX2_X2 U16067 ( .A(decode_regfile_intregs_20__22_), .B(
        decode_regfile_intregs_21__22_), .S(n12945), .Z(n11629) );
  MUX2_X2 U16068 ( .A(n11629), .B(n11628), .S(n13037), .Z(n11630) );
  MUX2_X2 U16069 ( .A(decode_regfile_intregs_18__22_), .B(
        decode_regfile_intregs_19__22_), .S(n12945), .Z(n11631) );
  MUX2_X2 U16070 ( .A(decode_regfile_intregs_16__22_), .B(
        decode_regfile_intregs_17__22_), .S(n12945), .Z(n11632) );
  MUX2_X2 U16071 ( .A(n11632), .B(n11631), .S(n13037), .Z(n11633) );
  MUX2_X2 U16072 ( .A(n11633), .B(n11630), .S(n13069), .Z(n11634) );
  MUX2_X2 U16073 ( .A(n11634), .B(n11627), .S(n13087), .Z(n11635) );
  MUX2_X2 U16074 ( .A(decode_regfile_intregs_14__22_), .B(
        decode_regfile_intregs_15__22_), .S(n12945), .Z(n11636) );
  MUX2_X2 U16075 ( .A(decode_regfile_intregs_12__22_), .B(
        decode_regfile_intregs_13__22_), .S(n12945), .Z(n11637) );
  MUX2_X2 U16076 ( .A(n11637), .B(n11636), .S(n13037), .Z(n11638) );
  MUX2_X2 U16077 ( .A(decode_regfile_intregs_10__22_), .B(
        decode_regfile_intregs_11__22_), .S(n12945), .Z(n11639) );
  MUX2_X2 U16078 ( .A(decode_regfile_intregs_8__22_), .B(
        decode_regfile_intregs_9__22_), .S(n12945), .Z(n11640) );
  MUX2_X2 U16079 ( .A(n11640), .B(n11639), .S(n13037), .Z(n11641) );
  MUX2_X2 U16080 ( .A(n11641), .B(n11638), .S(n13069), .Z(n11642) );
  MUX2_X2 U16081 ( .A(decode_regfile_intregs_6__22_), .B(
        decode_regfile_intregs_7__22_), .S(n12946), .Z(n11643) );
  MUX2_X2 U16082 ( .A(decode_regfile_intregs_4__22_), .B(
        decode_regfile_intregs_5__22_), .S(n12946), .Z(n11644) );
  MUX2_X2 U16083 ( .A(n11644), .B(n11643), .S(n13038), .Z(n11645) );
  MUX2_X2 U16084 ( .A(decode_regfile_intregs_2__22_), .B(
        decode_regfile_intregs_3__22_), .S(n12946), .Z(n11646) );
  MUX2_X2 U16085 ( .A(decode_regfile_intregs_0__22_), .B(
        decode_regfile_intregs_1__22_), .S(n12946), .Z(n11647) );
  MUX2_X2 U16086 ( .A(n11647), .B(n11646), .S(n13038), .Z(n11648) );
  MUX2_X2 U16087 ( .A(n11648), .B(n11645), .S(n13070), .Z(n11649) );
  MUX2_X2 U16088 ( .A(n11649), .B(n11642), .S(n13087), .Z(n11650) );
  MUX2_X2 U16089 ( .A(n11650), .B(n11635), .S(n13098), .Z(decode_regfile_N109)
         );
  MUX2_X2 U16090 ( .A(decode_regfile_intregs_30__23_), .B(
        decode_regfile_intregs_31__23_), .S(n12946), .Z(n11651) );
  MUX2_X2 U16091 ( .A(decode_regfile_intregs_28__23_), .B(
        decode_regfile_intregs_29__23_), .S(n12946), .Z(n11652) );
  MUX2_X2 U16092 ( .A(n11652), .B(n11651), .S(n13038), .Z(n11653) );
  MUX2_X2 U16093 ( .A(decode_regfile_intregs_26__23_), .B(
        decode_regfile_intregs_27__23_), .S(n12946), .Z(n11654) );
  MUX2_X2 U16094 ( .A(decode_regfile_intregs_24__23_), .B(
        decode_regfile_intregs_25__23_), .S(n12946), .Z(n11655) );
  MUX2_X2 U16095 ( .A(n11655), .B(n11654), .S(n13038), .Z(n11656) );
  MUX2_X2 U16096 ( .A(n11656), .B(n11653), .S(n13070), .Z(n11657) );
  MUX2_X2 U16097 ( .A(decode_regfile_intregs_22__23_), .B(
        decode_regfile_intregs_23__23_), .S(n12946), .Z(n11658) );
  MUX2_X2 U16098 ( .A(decode_regfile_intregs_20__23_), .B(
        decode_regfile_intregs_21__23_), .S(n12946), .Z(n11659) );
  MUX2_X2 U16099 ( .A(n11659), .B(n11658), .S(n13038), .Z(n11660) );
  MUX2_X2 U16100 ( .A(decode_regfile_intregs_18__23_), .B(
        decode_regfile_intregs_19__23_), .S(n12946), .Z(n11661) );
  MUX2_X2 U16101 ( .A(decode_regfile_intregs_16__23_), .B(
        decode_regfile_intregs_17__23_), .S(n12947), .Z(n11662) );
  MUX2_X2 U16102 ( .A(n11662), .B(n11661), .S(n13038), .Z(n11663) );
  MUX2_X2 U16103 ( .A(n11663), .B(n11660), .S(n13070), .Z(n11664) );
  MUX2_X2 U16104 ( .A(n11664), .B(n11657), .S(n13087), .Z(n11665) );
  MUX2_X2 U16105 ( .A(decode_regfile_intregs_14__23_), .B(
        decode_regfile_intregs_15__23_), .S(n12947), .Z(n11666) );
  MUX2_X2 U16106 ( .A(decode_regfile_intregs_12__23_), .B(
        decode_regfile_intregs_13__23_), .S(n12947), .Z(n11667) );
  MUX2_X2 U16107 ( .A(n11667), .B(n11666), .S(n13038), .Z(n11668) );
  MUX2_X2 U16108 ( .A(decode_regfile_intregs_10__23_), .B(
        decode_regfile_intregs_11__23_), .S(n12947), .Z(n11669) );
  MUX2_X2 U16109 ( .A(decode_regfile_intregs_8__23_), .B(
        decode_regfile_intregs_9__23_), .S(n12947), .Z(n11670) );
  MUX2_X2 U16110 ( .A(n11670), .B(n11669), .S(n13038), .Z(n11671) );
  MUX2_X2 U16111 ( .A(n11671), .B(n11668), .S(n13070), .Z(n11672) );
  MUX2_X2 U16112 ( .A(decode_regfile_intregs_6__23_), .B(
        decode_regfile_intregs_7__23_), .S(n12947), .Z(n11673) );
  MUX2_X2 U16113 ( .A(decode_regfile_intregs_4__23_), .B(
        decode_regfile_intregs_5__23_), .S(n12947), .Z(n11674) );
  MUX2_X2 U16114 ( .A(n11674), .B(n11673), .S(n13038), .Z(n11675) );
  MUX2_X2 U16115 ( .A(decode_regfile_intregs_2__23_), .B(
        decode_regfile_intregs_3__23_), .S(n12947), .Z(n11676) );
  MUX2_X2 U16116 ( .A(decode_regfile_intregs_0__23_), .B(
        decode_regfile_intregs_1__23_), .S(n12947), .Z(n11677) );
  MUX2_X2 U16117 ( .A(n11677), .B(n11676), .S(n13038), .Z(n11678) );
  MUX2_X2 U16118 ( .A(n11678), .B(n11675), .S(n13070), .Z(n11679) );
  MUX2_X2 U16119 ( .A(n11679), .B(n11672), .S(n13087), .Z(n11680) );
  MUX2_X2 U16120 ( .A(n11680), .B(n11665), .S(n13098), .Z(decode_regfile_N108)
         );
  MUX2_X2 U16121 ( .A(decode_regfile_intregs_30__24_), .B(
        decode_regfile_intregs_31__24_), .S(n12947), .Z(n11681) );
  MUX2_X2 U16122 ( .A(decode_regfile_intregs_28__24_), .B(
        decode_regfile_intregs_29__24_), .S(n12947), .Z(n11682) );
  MUX2_X2 U16123 ( .A(n11682), .B(n11681), .S(n13038), .Z(n11683) );
  MUX2_X2 U16124 ( .A(decode_regfile_intregs_26__24_), .B(
        decode_regfile_intregs_27__24_), .S(n12948), .Z(n11684) );
  MUX2_X2 U16125 ( .A(decode_regfile_intregs_24__24_), .B(
        decode_regfile_intregs_25__24_), .S(n12948), .Z(n11685) );
  MUX2_X2 U16126 ( .A(n11685), .B(n11684), .S(n13039), .Z(n11686) );
  MUX2_X2 U16127 ( .A(n11686), .B(n11683), .S(n13070), .Z(n11687) );
  MUX2_X2 U16128 ( .A(decode_regfile_intregs_22__24_), .B(
        decode_regfile_intregs_23__24_), .S(n12948), .Z(n11688) );
  MUX2_X2 U16129 ( .A(decode_regfile_intregs_20__24_), .B(
        decode_regfile_intregs_21__24_), .S(n12948), .Z(n11689) );
  MUX2_X2 U16130 ( .A(n11689), .B(n11688), .S(n13039), .Z(n11690) );
  MUX2_X2 U16131 ( .A(decode_regfile_intregs_18__24_), .B(
        decode_regfile_intregs_19__24_), .S(n12948), .Z(n11691) );
  MUX2_X2 U16132 ( .A(decode_regfile_intregs_16__24_), .B(
        decode_regfile_intregs_17__24_), .S(n12948), .Z(n11692) );
  MUX2_X2 U16133 ( .A(n11692), .B(n11691), .S(n13039), .Z(n11693) );
  MUX2_X2 U16134 ( .A(n11693), .B(n11690), .S(n13070), .Z(n11694) );
  MUX2_X2 U16135 ( .A(n11694), .B(n11687), .S(n13087), .Z(n11695) );
  MUX2_X2 U16136 ( .A(decode_regfile_intregs_14__24_), .B(
        decode_regfile_intregs_15__24_), .S(n12948), .Z(n11696) );
  MUX2_X2 U16137 ( .A(decode_regfile_intregs_12__24_), .B(
        decode_regfile_intregs_13__24_), .S(n12948), .Z(n11697) );
  MUX2_X2 U16138 ( .A(n11697), .B(n11696), .S(n13039), .Z(n11698) );
  MUX2_X2 U16139 ( .A(decode_regfile_intregs_10__24_), .B(
        decode_regfile_intregs_11__24_), .S(n12948), .Z(n11699) );
  MUX2_X2 U16140 ( .A(decode_regfile_intregs_8__24_), .B(
        decode_regfile_intregs_9__24_), .S(n12948), .Z(n11700) );
  MUX2_X2 U16141 ( .A(n11700), .B(n11699), .S(n13039), .Z(n11701) );
  MUX2_X2 U16142 ( .A(n11701), .B(n11698), .S(n13070), .Z(n11702) );
  MUX2_X2 U16143 ( .A(decode_regfile_intregs_6__24_), .B(
        decode_regfile_intregs_7__24_), .S(n12948), .Z(n11703) );
  MUX2_X2 U16144 ( .A(decode_regfile_intregs_4__24_), .B(
        decode_regfile_intregs_5__24_), .S(n12949), .Z(n11704) );
  MUX2_X2 U16145 ( .A(n11704), .B(n11703), .S(n13039), .Z(n11705) );
  MUX2_X2 U16146 ( .A(decode_regfile_intregs_2__24_), .B(
        decode_regfile_intregs_3__24_), .S(n12949), .Z(n11706) );
  MUX2_X2 U16147 ( .A(decode_regfile_intregs_0__24_), .B(
        decode_regfile_intregs_1__24_), .S(n12949), .Z(n11707) );
  MUX2_X2 U16148 ( .A(n11707), .B(n11706), .S(n13039), .Z(n11708) );
  MUX2_X2 U16149 ( .A(n11708), .B(n11705), .S(n13070), .Z(n11709) );
  MUX2_X2 U16150 ( .A(n11709), .B(n11702), .S(n13087), .Z(n11710) );
  MUX2_X2 U16151 ( .A(n11710), .B(n11695), .S(n13098), .Z(decode_regfile_N107)
         );
  MUX2_X2 U16152 ( .A(decode_regfile_intregs_30__25_), .B(
        decode_regfile_intregs_31__25_), .S(n12949), .Z(n11711) );
  MUX2_X2 U16153 ( .A(decode_regfile_intregs_28__25_), .B(
        decode_regfile_intregs_29__25_), .S(n12949), .Z(n11712) );
  MUX2_X2 U16154 ( .A(n11712), .B(n11711), .S(n13039), .Z(n11713) );
  MUX2_X2 U16155 ( .A(decode_regfile_intregs_26__25_), .B(
        decode_regfile_intregs_27__25_), .S(n12949), .Z(n11714) );
  MUX2_X2 U16156 ( .A(decode_regfile_intregs_24__25_), .B(
        decode_regfile_intregs_25__25_), .S(n12949), .Z(n11715) );
  MUX2_X2 U16157 ( .A(n11715), .B(n11714), .S(n13039), .Z(n11716) );
  MUX2_X2 U16158 ( .A(n11716), .B(n11713), .S(n13070), .Z(n11717) );
  MUX2_X2 U16159 ( .A(decode_regfile_intregs_22__25_), .B(
        decode_regfile_intregs_23__25_), .S(n12949), .Z(n11718) );
  MUX2_X2 U16160 ( .A(decode_regfile_intregs_20__25_), .B(
        decode_regfile_intregs_21__25_), .S(n12949), .Z(n11719) );
  MUX2_X2 U16161 ( .A(n11719), .B(n11718), .S(n13039), .Z(n11720) );
  MUX2_X2 U16162 ( .A(decode_regfile_intregs_18__25_), .B(
        decode_regfile_intregs_19__25_), .S(n12949), .Z(n11721) );
  MUX2_X2 U16163 ( .A(decode_regfile_intregs_16__25_), .B(
        decode_regfile_intregs_17__25_), .S(n12949), .Z(n11722) );
  MUX2_X2 U16164 ( .A(n11722), .B(n11721), .S(n13039), .Z(n11723) );
  MUX2_X2 U16165 ( .A(n11723), .B(n11720), .S(n13070), .Z(n11724) );
  MUX2_X2 U16166 ( .A(n11724), .B(n11717), .S(n13087), .Z(n11725) );
  MUX2_X2 U16167 ( .A(decode_regfile_intregs_14__25_), .B(
        decode_regfile_intregs_15__25_), .S(n12950), .Z(n11726) );
  MUX2_X2 U16168 ( .A(decode_regfile_intregs_12__25_), .B(
        decode_regfile_intregs_13__25_), .S(n12950), .Z(n11727) );
  MUX2_X2 U16169 ( .A(n11727), .B(n11726), .S(n13040), .Z(n11728) );
  MUX2_X2 U16170 ( .A(decode_regfile_intregs_10__25_), .B(
        decode_regfile_intregs_11__25_), .S(n12950), .Z(n11729) );
  MUX2_X2 U16171 ( .A(decode_regfile_intregs_8__25_), .B(
        decode_regfile_intregs_9__25_), .S(n12950), .Z(n11730) );
  MUX2_X2 U16172 ( .A(n11730), .B(n11729), .S(n13040), .Z(n11731) );
  MUX2_X2 U16173 ( .A(n11731), .B(n11728), .S(n13071), .Z(n11732) );
  MUX2_X2 U16174 ( .A(decode_regfile_intregs_6__25_), .B(
        decode_regfile_intregs_7__25_), .S(n12950), .Z(n11733) );
  MUX2_X2 U16175 ( .A(decode_regfile_intregs_4__25_), .B(
        decode_regfile_intregs_5__25_), .S(n12950), .Z(n11734) );
  MUX2_X2 U16176 ( .A(n11734), .B(n11733), .S(n13040), .Z(n11735) );
  MUX2_X2 U16177 ( .A(decode_regfile_intregs_2__25_), .B(
        decode_regfile_intregs_3__25_), .S(n12950), .Z(n11736) );
  MUX2_X2 U16178 ( .A(decode_regfile_intregs_0__25_), .B(
        decode_regfile_intregs_1__25_), .S(n12950), .Z(n11737) );
  MUX2_X2 U16179 ( .A(n11737), .B(n11736), .S(n13040), .Z(n11738) );
  MUX2_X2 U16180 ( .A(n11738), .B(n11735), .S(n13071), .Z(n11739) );
  MUX2_X2 U16181 ( .A(n11739), .B(n11732), .S(n13088), .Z(n11740) );
  MUX2_X2 U16182 ( .A(n11740), .B(n11725), .S(n13098), .Z(decode_regfile_N106)
         );
  MUX2_X2 U16183 ( .A(decode_regfile_intregs_30__26_), .B(
        decode_regfile_intregs_31__26_), .S(n12950), .Z(n11741) );
  MUX2_X2 U16184 ( .A(decode_regfile_intregs_28__26_), .B(
        decode_regfile_intregs_29__26_), .S(n12950), .Z(n11742) );
  MUX2_X2 U16185 ( .A(n11742), .B(n11741), .S(n13040), .Z(n11743) );
  MUX2_X2 U16186 ( .A(decode_regfile_intregs_26__26_), .B(
        decode_regfile_intregs_27__26_), .S(n12950), .Z(n11744) );
  MUX2_X2 U16187 ( .A(decode_regfile_intregs_24__26_), .B(
        decode_regfile_intregs_25__26_), .S(n12951), .Z(n11745) );
  MUX2_X2 U16188 ( .A(n11745), .B(n11744), .S(n13040), .Z(n11746) );
  MUX2_X2 U16189 ( .A(n11746), .B(n11743), .S(n13071), .Z(n11747) );
  MUX2_X2 U16190 ( .A(decode_regfile_intregs_22__26_), .B(
        decode_regfile_intregs_23__26_), .S(n12951), .Z(n11748) );
  MUX2_X2 U16191 ( .A(decode_regfile_intregs_20__26_), .B(
        decode_regfile_intregs_21__26_), .S(n12951), .Z(n11749) );
  MUX2_X2 U16192 ( .A(n11749), .B(n11748), .S(n13040), .Z(n11750) );
  MUX2_X2 U16193 ( .A(decode_regfile_intregs_18__26_), .B(
        decode_regfile_intregs_19__26_), .S(n12951), .Z(n11751) );
  MUX2_X2 U16194 ( .A(decode_regfile_intregs_16__26_), .B(
        decode_regfile_intregs_17__26_), .S(n12951), .Z(n11752) );
  MUX2_X2 U16195 ( .A(n11752), .B(n11751), .S(n13040), .Z(n11753) );
  MUX2_X2 U16196 ( .A(n11753), .B(n11750), .S(n13071), .Z(n11754) );
  MUX2_X2 U16197 ( .A(n11754), .B(n11747), .S(n13088), .Z(n11755) );
  MUX2_X2 U16198 ( .A(decode_regfile_intregs_14__26_), .B(
        decode_regfile_intregs_15__26_), .S(n12951), .Z(n11756) );
  MUX2_X2 U16199 ( .A(decode_regfile_intregs_12__26_), .B(
        decode_regfile_intregs_13__26_), .S(n12951), .Z(n11757) );
  MUX2_X2 U16200 ( .A(n11757), .B(n11756), .S(n13040), .Z(n11758) );
  MUX2_X2 U16201 ( .A(decode_regfile_intregs_10__26_), .B(
        decode_regfile_intregs_11__26_), .S(n12951), .Z(n11759) );
  MUX2_X2 U16202 ( .A(decode_regfile_intregs_8__26_), .B(
        decode_regfile_intregs_9__26_), .S(n12951), .Z(n11760) );
  MUX2_X2 U16203 ( .A(n11760), .B(n11759), .S(n13040), .Z(n11761) );
  MUX2_X2 U16204 ( .A(n11761), .B(n11758), .S(n13071), .Z(n11762) );
  MUX2_X2 U16205 ( .A(decode_regfile_intregs_6__26_), .B(
        decode_regfile_intregs_7__26_), .S(n12951), .Z(n11763) );
  MUX2_X2 U16206 ( .A(decode_regfile_intregs_4__26_), .B(
        decode_regfile_intregs_5__26_), .S(n12951), .Z(n11764) );
  MUX2_X2 U16207 ( .A(n11764), .B(n11763), .S(n13040), .Z(n11765) );
  MUX2_X2 U16208 ( .A(decode_regfile_intregs_2__26_), .B(
        decode_regfile_intregs_3__26_), .S(n12952), .Z(n11766) );
  MUX2_X2 U16209 ( .A(decode_regfile_intregs_0__26_), .B(
        decode_regfile_intregs_1__26_), .S(n12952), .Z(n11767) );
  MUX2_X2 U16210 ( .A(n11767), .B(n11766), .S(n13041), .Z(n11768) );
  MUX2_X2 U16211 ( .A(n11768), .B(n11765), .S(n13071), .Z(n11769) );
  MUX2_X2 U16212 ( .A(n11769), .B(n11762), .S(n13088), .Z(n11770) );
  MUX2_X2 U16213 ( .A(n11770), .B(n11755), .S(n13098), .Z(decode_regfile_N105)
         );
  MUX2_X2 U16214 ( .A(decode_regfile_intregs_30__27_), .B(
        decode_regfile_intregs_31__27_), .S(n12952), .Z(n11771) );
  MUX2_X2 U16215 ( .A(decode_regfile_intregs_28__27_), .B(
        decode_regfile_intregs_29__27_), .S(n12952), .Z(n11772) );
  MUX2_X2 U16216 ( .A(n11772), .B(n11771), .S(n13041), .Z(n11773) );
  MUX2_X2 U16217 ( .A(decode_regfile_intregs_26__27_), .B(
        decode_regfile_intregs_27__27_), .S(n12952), .Z(n11774) );
  MUX2_X2 U16218 ( .A(decode_regfile_intregs_24__27_), .B(
        decode_regfile_intregs_25__27_), .S(n12952), .Z(n11775) );
  MUX2_X2 U16219 ( .A(n11775), .B(n11774), .S(n13041), .Z(n11776) );
  MUX2_X2 U16220 ( .A(n11776), .B(n11773), .S(n13071), .Z(n11777) );
  MUX2_X2 U16221 ( .A(decode_regfile_intregs_22__27_), .B(
        decode_regfile_intregs_23__27_), .S(n12952), .Z(n11778) );
  MUX2_X2 U16222 ( .A(decode_regfile_intregs_20__27_), .B(
        decode_regfile_intregs_21__27_), .S(n12952), .Z(n11779) );
  MUX2_X2 U16223 ( .A(n11779), .B(n11778), .S(n13041), .Z(n11780) );
  MUX2_X2 U16224 ( .A(decode_regfile_intregs_18__27_), .B(
        decode_regfile_intregs_19__27_), .S(n12952), .Z(n11781) );
  MUX2_X2 U16225 ( .A(decode_regfile_intregs_16__27_), .B(
        decode_regfile_intregs_17__27_), .S(n12952), .Z(n11782) );
  MUX2_X2 U16226 ( .A(n11782), .B(n11781), .S(n13041), .Z(n11783) );
  MUX2_X2 U16227 ( .A(n11783), .B(n11780), .S(n13071), .Z(n11784) );
  MUX2_X2 U16228 ( .A(n11784), .B(n11777), .S(n13088), .Z(n11785) );
  MUX2_X2 U16229 ( .A(decode_regfile_intregs_14__27_), .B(
        decode_regfile_intregs_15__27_), .S(n12952), .Z(n11786) );
  MUX2_X2 U16230 ( .A(decode_regfile_intregs_12__27_), .B(
        decode_regfile_intregs_13__27_), .S(n12953), .Z(n11787) );
  MUX2_X2 U16231 ( .A(n11787), .B(n11786), .S(n13041), .Z(n11788) );
  MUX2_X2 U16232 ( .A(decode_regfile_intregs_10__27_), .B(
        decode_regfile_intregs_11__27_), .S(n12953), .Z(n11789) );
  MUX2_X2 U16233 ( .A(decode_regfile_intregs_8__27_), .B(
        decode_regfile_intregs_9__27_), .S(n12953), .Z(n11790) );
  MUX2_X2 U16234 ( .A(n11790), .B(n11789), .S(n13041), .Z(n11791) );
  MUX2_X2 U16235 ( .A(n11791), .B(n11788), .S(n13071), .Z(n11792) );
  MUX2_X2 U16236 ( .A(decode_regfile_intregs_6__27_), .B(
        decode_regfile_intregs_7__27_), .S(n12953), .Z(n11793) );
  MUX2_X2 U16237 ( .A(decode_regfile_intregs_4__27_), .B(
        decode_regfile_intregs_5__27_), .S(n12953), .Z(n11794) );
  MUX2_X2 U16238 ( .A(n11794), .B(n11793), .S(n13041), .Z(n11795) );
  MUX2_X2 U16239 ( .A(decode_regfile_intregs_2__27_), .B(
        decode_regfile_intregs_3__27_), .S(n12953), .Z(n11796) );
  MUX2_X2 U16240 ( .A(decode_regfile_intregs_0__27_), .B(
        decode_regfile_intregs_1__27_), .S(n12953), .Z(n11797) );
  MUX2_X2 U16241 ( .A(n11797), .B(n11796), .S(n13041), .Z(n11798) );
  MUX2_X2 U16242 ( .A(n11798), .B(n11795), .S(n13071), .Z(n11799) );
  MUX2_X2 U16243 ( .A(n11799), .B(n11792), .S(n13088), .Z(n11800) );
  MUX2_X2 U16244 ( .A(n11800), .B(n11785), .S(n13098), .Z(decode_regfile_N104)
         );
  MUX2_X2 U16245 ( .A(decode_regfile_intregs_30__28_), .B(
        decode_regfile_intregs_31__28_), .S(n12953), .Z(n11801) );
  MUX2_X2 U16246 ( .A(decode_regfile_intregs_28__28_), .B(
        decode_regfile_intregs_29__28_), .S(n12953), .Z(n11802) );
  MUX2_X2 U16247 ( .A(n11802), .B(n11801), .S(n13041), .Z(n11803) );
  MUX2_X2 U16248 ( .A(decode_regfile_intregs_26__28_), .B(
        decode_regfile_intregs_27__28_), .S(n12953), .Z(n11804) );
  MUX2_X2 U16249 ( .A(decode_regfile_intregs_24__28_), .B(
        decode_regfile_intregs_25__28_), .S(n12953), .Z(n11805) );
  MUX2_X2 U16250 ( .A(n11805), .B(n11804), .S(n13041), .Z(n11806) );
  MUX2_X2 U16251 ( .A(n11806), .B(n11803), .S(n13071), .Z(n11807) );
  MUX2_X2 U16252 ( .A(decode_regfile_intregs_22__28_), .B(
        decode_regfile_intregs_23__28_), .S(n12954), .Z(n11808) );
  MUX2_X2 U16253 ( .A(decode_regfile_intregs_20__28_), .B(
        decode_regfile_intregs_21__28_), .S(n12954), .Z(n11809) );
  MUX2_X2 U16254 ( .A(n11809), .B(n11808), .S(n13042), .Z(n11810) );
  MUX2_X2 U16255 ( .A(decode_regfile_intregs_18__28_), .B(
        decode_regfile_intregs_19__28_), .S(n12954), .Z(n11811) );
  MUX2_X2 U16256 ( .A(decode_regfile_intregs_16__28_), .B(
        decode_regfile_intregs_17__28_), .S(n12954), .Z(n11812) );
  MUX2_X2 U16257 ( .A(n11812), .B(n11811), .S(n13042), .Z(n11813) );
  MUX2_X2 U16258 ( .A(n11813), .B(n11810), .S(n13072), .Z(n11814) );
  MUX2_X2 U16259 ( .A(n11814), .B(n11807), .S(n13088), .Z(n11815) );
  MUX2_X2 U16260 ( .A(decode_regfile_intregs_14__28_), .B(
        decode_regfile_intregs_15__28_), .S(n12954), .Z(n11816) );
  MUX2_X2 U16261 ( .A(decode_regfile_intregs_12__28_), .B(
        decode_regfile_intregs_13__28_), .S(n12954), .Z(n11817) );
  MUX2_X2 U16262 ( .A(n11817), .B(n11816), .S(n13042), .Z(n11818) );
  MUX2_X2 U16263 ( .A(decode_regfile_intregs_10__28_), .B(
        decode_regfile_intregs_11__28_), .S(n12954), .Z(n11819) );
  MUX2_X2 U16264 ( .A(decode_regfile_intregs_8__28_), .B(
        decode_regfile_intregs_9__28_), .S(n12954), .Z(n11820) );
  MUX2_X2 U16265 ( .A(n11820), .B(n11819), .S(n13042), .Z(n11821) );
  MUX2_X2 U16266 ( .A(n11821), .B(n11818), .S(n13072), .Z(n11822) );
  MUX2_X2 U16267 ( .A(decode_regfile_intregs_6__28_), .B(
        decode_regfile_intregs_7__28_), .S(n12954), .Z(n11823) );
  MUX2_X2 U16268 ( .A(decode_regfile_intregs_4__28_), .B(
        decode_regfile_intregs_5__28_), .S(n12954), .Z(n11824) );
  MUX2_X2 U16269 ( .A(n11824), .B(n11823), .S(n13042), .Z(n11825) );
  MUX2_X2 U16270 ( .A(decode_regfile_intregs_2__28_), .B(
        decode_regfile_intregs_3__28_), .S(n12954), .Z(n11826) );
  MUX2_X2 U16271 ( .A(decode_regfile_intregs_0__28_), .B(
        decode_regfile_intregs_1__28_), .S(n12955), .Z(n11827) );
  MUX2_X2 U16272 ( .A(n11827), .B(n11826), .S(n13042), .Z(n11828) );
  MUX2_X2 U16273 ( .A(n11828), .B(n11825), .S(n13072), .Z(n11829) );
  MUX2_X2 U16274 ( .A(n11829), .B(n11822), .S(n13088), .Z(n11830) );
  MUX2_X2 U16275 ( .A(n11830), .B(n11815), .S(n13098), .Z(decode_regfile_N103)
         );
  MUX2_X2 U16276 ( .A(decode_regfile_intregs_30__29_), .B(
        decode_regfile_intregs_31__29_), .S(n12955), .Z(n11831) );
  MUX2_X2 U16277 ( .A(decode_regfile_intregs_28__29_), .B(
        decode_regfile_intregs_29__29_), .S(n12955), .Z(n11832) );
  MUX2_X2 U16278 ( .A(n11832), .B(n11831), .S(n13042), .Z(n11833) );
  MUX2_X2 U16279 ( .A(decode_regfile_intregs_26__29_), .B(
        decode_regfile_intregs_27__29_), .S(n12955), .Z(n11834) );
  MUX2_X2 U16280 ( .A(decode_regfile_intregs_24__29_), .B(
        decode_regfile_intregs_25__29_), .S(n12955), .Z(n11835) );
  MUX2_X2 U16281 ( .A(n11835), .B(n11834), .S(n13042), .Z(n11836) );
  MUX2_X2 U16282 ( .A(n11836), .B(n11833), .S(n13072), .Z(n11837) );
  MUX2_X2 U16283 ( .A(decode_regfile_intregs_22__29_), .B(
        decode_regfile_intregs_23__29_), .S(n12955), .Z(n11838) );
  MUX2_X2 U16284 ( .A(decode_regfile_intregs_20__29_), .B(
        decode_regfile_intregs_21__29_), .S(n12955), .Z(n11839) );
  MUX2_X2 U16285 ( .A(n11839), .B(n11838), .S(n13042), .Z(n11840) );
  MUX2_X2 U16286 ( .A(decode_regfile_intregs_18__29_), .B(
        decode_regfile_intregs_19__29_), .S(n12955), .Z(n11841) );
  MUX2_X2 U16287 ( .A(decode_regfile_intregs_16__29_), .B(
        decode_regfile_intregs_17__29_), .S(n12955), .Z(n11842) );
  MUX2_X2 U16288 ( .A(n11842), .B(n11841), .S(n13042), .Z(n11843) );
  MUX2_X2 U16289 ( .A(n11843), .B(n11840), .S(n13072), .Z(n11844) );
  MUX2_X2 U16290 ( .A(n11844), .B(n11837), .S(n13088), .Z(n11845) );
  MUX2_X2 U16291 ( .A(decode_regfile_intregs_14__29_), .B(
        decode_regfile_intregs_15__29_), .S(n12955), .Z(n11846) );
  MUX2_X2 U16292 ( .A(decode_regfile_intregs_12__29_), .B(
        decode_regfile_intregs_13__29_), .S(n12955), .Z(n11847) );
  MUX2_X2 U16293 ( .A(n11847), .B(n11846), .S(n13042), .Z(n11848) );
  MUX2_X2 U16294 ( .A(decode_regfile_intregs_10__29_), .B(
        decode_regfile_intregs_11__29_), .S(n12956), .Z(n11849) );
  MUX2_X2 U16295 ( .A(decode_regfile_intregs_8__29_), .B(
        decode_regfile_intregs_9__29_), .S(n12956), .Z(n11850) );
  MUX2_X2 U16296 ( .A(n11850), .B(n11849), .S(n13043), .Z(n11851) );
  MUX2_X2 U16297 ( .A(n11851), .B(n11848), .S(n13072), .Z(n11852) );
  MUX2_X2 U16298 ( .A(decode_regfile_intregs_6__29_), .B(
        decode_regfile_intregs_7__29_), .S(n12956), .Z(n11853) );
  MUX2_X2 U16299 ( .A(decode_regfile_intregs_4__29_), .B(
        decode_regfile_intregs_5__29_), .S(n12956), .Z(n11854) );
  MUX2_X2 U16300 ( .A(n11854), .B(n11853), .S(n13043), .Z(n11855) );
  MUX2_X2 U16301 ( .A(decode_regfile_intregs_2__29_), .B(
        decode_regfile_intregs_3__29_), .S(n12956), .Z(n11856) );
  MUX2_X2 U16302 ( .A(decode_regfile_intregs_0__29_), .B(
        decode_regfile_intregs_1__29_), .S(n12956), .Z(n11857) );
  MUX2_X2 U16303 ( .A(n11857), .B(n11856), .S(n13043), .Z(n11858) );
  MUX2_X2 U16304 ( .A(n11858), .B(n11855), .S(n13072), .Z(n11859) );
  MUX2_X2 U16305 ( .A(n11859), .B(n11852), .S(n13088), .Z(n11860) );
  MUX2_X2 U16306 ( .A(n11860), .B(n11845), .S(n13098), .Z(decode_regfile_N102)
         );
  MUX2_X2 U16307 ( .A(decode_regfile_intregs_30__30_), .B(
        decode_regfile_intregs_31__30_), .S(n12956), .Z(n11861) );
  MUX2_X2 U16308 ( .A(decode_regfile_intregs_28__30_), .B(
        decode_regfile_intregs_29__30_), .S(n12956), .Z(n11862) );
  MUX2_X2 U16309 ( .A(n11862), .B(n11861), .S(n13043), .Z(n11863) );
  MUX2_X2 U16310 ( .A(decode_regfile_intregs_26__30_), .B(
        decode_regfile_intregs_27__30_), .S(n12956), .Z(n11864) );
  MUX2_X2 U16311 ( .A(decode_regfile_intregs_24__30_), .B(
        decode_regfile_intregs_25__30_), .S(n12956), .Z(n11865) );
  MUX2_X2 U16312 ( .A(n11865), .B(n11864), .S(n13043), .Z(n11866) );
  MUX2_X2 U16313 ( .A(n11866), .B(n11863), .S(n13072), .Z(n11867) );
  MUX2_X2 U16314 ( .A(decode_regfile_intregs_22__30_), .B(
        decode_regfile_intregs_23__30_), .S(n12956), .Z(n11868) );
  MUX2_X2 U16315 ( .A(decode_regfile_intregs_20__30_), .B(
        decode_regfile_intregs_21__30_), .S(n12957), .Z(n11869) );
  MUX2_X2 U16316 ( .A(n11869), .B(n11868), .S(n13043), .Z(n11870) );
  MUX2_X2 U16317 ( .A(decode_regfile_intregs_18__30_), .B(
        decode_regfile_intregs_19__30_), .S(n12957), .Z(n11871) );
  MUX2_X2 U16318 ( .A(decode_regfile_intregs_16__30_), .B(
        decode_regfile_intregs_17__30_), .S(n12957), .Z(n11872) );
  MUX2_X2 U16319 ( .A(n11872), .B(n11871), .S(n13043), .Z(n11873) );
  MUX2_X2 U16320 ( .A(n11873), .B(n11870), .S(n13072), .Z(n11874) );
  MUX2_X2 U16321 ( .A(n11874), .B(n11867), .S(n13088), .Z(n11875) );
  MUX2_X2 U16322 ( .A(decode_regfile_intregs_14__30_), .B(
        decode_regfile_intregs_15__30_), .S(n12957), .Z(n11876) );
  MUX2_X2 U16323 ( .A(decode_regfile_intregs_12__30_), .B(
        decode_regfile_intregs_13__30_), .S(n12957), .Z(n11877) );
  MUX2_X2 U16324 ( .A(n11877), .B(n11876), .S(n13043), .Z(n11878) );
  MUX2_X2 U16325 ( .A(decode_regfile_intregs_10__30_), .B(
        decode_regfile_intregs_11__30_), .S(n12957), .Z(n11879) );
  MUX2_X2 U16326 ( .A(decode_regfile_intregs_8__30_), .B(
        decode_regfile_intregs_9__30_), .S(n12957), .Z(n11880) );
  MUX2_X2 U16327 ( .A(n11880), .B(n11879), .S(n13043), .Z(n11881) );
  MUX2_X2 U16328 ( .A(n11881), .B(n11878), .S(n13072), .Z(n11882) );
  MUX2_X2 U16329 ( .A(decode_regfile_intregs_6__30_), .B(
        decode_regfile_intregs_7__30_), .S(n12957), .Z(n11883) );
  MUX2_X2 U16330 ( .A(decode_regfile_intregs_4__30_), .B(
        decode_regfile_intregs_5__30_), .S(n12957), .Z(n11884) );
  MUX2_X2 U16331 ( .A(n11884), .B(n11883), .S(n13043), .Z(n11885) );
  MUX2_X2 U16332 ( .A(decode_regfile_intregs_2__30_), .B(
        decode_regfile_intregs_3__30_), .S(n12957), .Z(n11886) );
  MUX2_X2 U16333 ( .A(decode_regfile_intregs_0__30_), .B(
        decode_regfile_intregs_1__30_), .S(n12957), .Z(n11887) );
  MUX2_X2 U16334 ( .A(n11887), .B(n11886), .S(n13043), .Z(n11888) );
  MUX2_X2 U16335 ( .A(n11888), .B(n11885), .S(n13072), .Z(n11889) );
  MUX2_X2 U16336 ( .A(n11889), .B(n11882), .S(n13088), .Z(n11890) );
  MUX2_X2 U16337 ( .A(n11890), .B(n11875), .S(n13098), .Z(decode_regfile_N101)
         );
  MUX2_X2 U16338 ( .A(decode_regfile_intregs_30__31_), .B(
        decode_regfile_intregs_31__31_), .S(n12958), .Z(n11891) );
  MUX2_X2 U16339 ( .A(decode_regfile_intregs_28__31_), .B(
        decode_regfile_intregs_29__31_), .S(n12958), .Z(n11892) );
  MUX2_X2 U16340 ( .A(n11892), .B(n11891), .S(n13013), .Z(n11893) );
  MUX2_X2 U16341 ( .A(decode_regfile_intregs_26__31_), .B(
        decode_regfile_intregs_27__31_), .S(n12958), .Z(n11894) );
  MUX2_X2 U16342 ( .A(decode_regfile_intregs_24__31_), .B(
        decode_regfile_intregs_25__31_), .S(n12958), .Z(n11895) );
  MUX2_X2 U16343 ( .A(n11895), .B(n11894), .S(n13007), .Z(n11896) );
  MUX2_X2 U16344 ( .A(n11896), .B(n11893), .S(n13073), .Z(n11897) );
  MUX2_X2 U16345 ( .A(decode_regfile_intregs_22__31_), .B(
        decode_regfile_intregs_23__31_), .S(n12958), .Z(n11898) );
  MUX2_X2 U16346 ( .A(decode_regfile_intregs_20__31_), .B(
        decode_regfile_intregs_21__31_), .S(n12958), .Z(n11899) );
  MUX2_X2 U16347 ( .A(n11899), .B(n11898), .S(n13020), .Z(n11900) );
  MUX2_X2 U16348 ( .A(decode_regfile_intregs_18__31_), .B(
        decode_regfile_intregs_19__31_), .S(n12958), .Z(n11901) );
  MUX2_X2 U16349 ( .A(decode_regfile_intregs_16__31_), .B(
        decode_regfile_intregs_17__31_), .S(n12958), .Z(n11902) );
  MUX2_X2 U16350 ( .A(n11902), .B(n11901), .S(n13018), .Z(n11903) );
  MUX2_X2 U16351 ( .A(n11903), .B(n11900), .S(n13073), .Z(n11904) );
  MUX2_X2 U16352 ( .A(n11904), .B(n11897), .S(n13089), .Z(n11905) );
  MUX2_X2 U16353 ( .A(decode_regfile_intregs_14__31_), .B(
        decode_regfile_intregs_15__31_), .S(n12958), .Z(n11906) );
  MUX2_X2 U16354 ( .A(decode_regfile_intregs_12__31_), .B(
        decode_regfile_intregs_13__31_), .S(n12958), .Z(n11907) );
  MUX2_X2 U16355 ( .A(n11907), .B(n11906), .S(n13016), .Z(n11908) );
  MUX2_X2 U16356 ( .A(decode_regfile_intregs_10__31_), .B(
        decode_regfile_intregs_11__31_), .S(n12958), .Z(n11909) );
  MUX2_X2 U16357 ( .A(decode_regfile_intregs_8__31_), .B(
        decode_regfile_intregs_9__31_), .S(n12959), .Z(n11910) );
  MUX2_X2 U16358 ( .A(n11910), .B(n11909), .S(n13015), .Z(n11911) );
  MUX2_X2 U16359 ( .A(n11911), .B(n11908), .S(n13073), .Z(n11912) );
  MUX2_X2 U16360 ( .A(decode_regfile_intregs_6__31_), .B(
        decode_regfile_intregs_7__31_), .S(n12959), .Z(n11913) );
  MUX2_X2 U16361 ( .A(decode_regfile_intregs_4__31_), .B(
        decode_regfile_intregs_5__31_), .S(n12959), .Z(n11914) );
  MUX2_X2 U16362 ( .A(n11914), .B(n11913), .S(n13009), .Z(n11915) );
  MUX2_X2 U16363 ( .A(decode_regfile_intregs_2__31_), .B(
        decode_regfile_intregs_3__31_), .S(n12959), .Z(n11916) );
  MUX2_X2 U16364 ( .A(decode_regfile_intregs_0__31_), .B(
        decode_regfile_intregs_1__31_), .S(n12959), .Z(n11917) );
  MUX2_X2 U16365 ( .A(n11917), .B(n11916), .S(n13012), .Z(n11918) );
  MUX2_X2 U16366 ( .A(n11918), .B(n11915), .S(n13073), .Z(n11919) );
  MUX2_X2 U16367 ( .A(n11919), .B(n11912), .S(n13089), .Z(n11920) );
  MUX2_X2 U16368 ( .A(n11920), .B(n11905), .S(n13099), .Z(decode_regfile_N100)
         );
  MUX2_X2 U16369 ( .A(decode_regfile_fpregs_30__0_), .B(
        decode_regfile_fpregs_31__0_), .S(n12959), .Z(n11921) );
  MUX2_X2 U16370 ( .A(decode_regfile_fpregs_28__0_), .B(
        decode_regfile_fpregs_29__0_), .S(n12959), .Z(n11922) );
  MUX2_X2 U16371 ( .A(n11922), .B(n11921), .S(n13014), .Z(n11923) );
  MUX2_X2 U16372 ( .A(decode_regfile_fpregs_26__0_), .B(
        decode_regfile_fpregs_27__0_), .S(n12959), .Z(n11924) );
  MUX2_X2 U16373 ( .A(decode_regfile_fpregs_24__0_), .B(
        decode_regfile_fpregs_25__0_), .S(n12959), .Z(n11925) );
  MUX2_X2 U16374 ( .A(n11925), .B(n11924), .S(n13019), .Z(n11926) );
  MUX2_X2 U16375 ( .A(n11926), .B(n11923), .S(n13073), .Z(n11927) );
  MUX2_X2 U16376 ( .A(decode_regfile_fpregs_22__0_), .B(
        decode_regfile_fpregs_23__0_), .S(n12959), .Z(n11928) );
  MUX2_X2 U16377 ( .A(decode_regfile_fpregs_20__0_), .B(
        decode_regfile_fpregs_21__0_), .S(n12959), .Z(n11929) );
  MUX2_X2 U16378 ( .A(n11929), .B(n11928), .S(n13017), .Z(n11930) );
  MUX2_X2 U16379 ( .A(decode_regfile_fpregs_18__0_), .B(
        decode_regfile_fpregs_19__0_), .S(n12960), .Z(n11931) );
  MUX2_X2 U16380 ( .A(decode_regfile_fpregs_16__0_), .B(
        decode_regfile_fpregs_17__0_), .S(n12960), .Z(n11932) );
  MUX2_X2 U16381 ( .A(n11932), .B(n11931), .S(n13044), .Z(n11933) );
  MUX2_X2 U16382 ( .A(n11933), .B(n11930), .S(n13073), .Z(n11934) );
  MUX2_X2 U16383 ( .A(n11934), .B(n11927), .S(n13089), .Z(n11935) );
  MUX2_X2 U16384 ( .A(decode_regfile_fpregs_14__0_), .B(
        decode_regfile_fpregs_15__0_), .S(n12960), .Z(n11936) );
  MUX2_X2 U16385 ( .A(decode_regfile_fpregs_12__0_), .B(
        decode_regfile_fpregs_13__0_), .S(n12960), .Z(n11937) );
  MUX2_X2 U16386 ( .A(n11937), .B(n11936), .S(n13044), .Z(n11938) );
  MUX2_X2 U16387 ( .A(decode_regfile_fpregs_10__0_), .B(
        decode_regfile_fpregs_11__0_), .S(n12960), .Z(n11939) );
  MUX2_X2 U16388 ( .A(decode_regfile_fpregs_8__0_), .B(
        decode_regfile_fpregs_9__0_), .S(n12960), .Z(n11940) );
  MUX2_X2 U16389 ( .A(n11940), .B(n11939), .S(n13044), .Z(n11941) );
  MUX2_X2 U16390 ( .A(n11941), .B(n11938), .S(n13073), .Z(n11942) );
  MUX2_X2 U16391 ( .A(decode_regfile_fpregs_6__0_), .B(
        decode_regfile_fpregs_7__0_), .S(n12960), .Z(n11943) );
  MUX2_X2 U16392 ( .A(decode_regfile_fpregs_4__0_), .B(
        decode_regfile_fpregs_5__0_), .S(n12960), .Z(n11944) );
  MUX2_X2 U16393 ( .A(n11944), .B(n11943), .S(n13044), .Z(n11945) );
  MUX2_X2 U16394 ( .A(decode_regfile_fpregs_2__0_), .B(
        decode_regfile_fpregs_3__0_), .S(n12960), .Z(n11946) );
  MUX2_X2 U16395 ( .A(decode_regfile_fpregs_0__0_), .B(
        decode_regfile_fpregs_1__0_), .S(n12960), .Z(n11947) );
  MUX2_X2 U16396 ( .A(n11947), .B(n11946), .S(n13044), .Z(n11948) );
  MUX2_X2 U16397 ( .A(n11948), .B(n11945), .S(n13073), .Z(n11949) );
  MUX2_X2 U16398 ( .A(n11949), .B(n11942), .S(n13089), .Z(n11950) );
  MUX2_X2 U16399 ( .A(n11950), .B(n11935), .S(n13099), .Z(decode_regfile_N163)
         );
  MUX2_X2 U16400 ( .A(decode_regfile_fpregs_30__1_), .B(
        decode_regfile_fpregs_31__1_), .S(n12960), .Z(n11951) );
  MUX2_X2 U16401 ( .A(decode_regfile_fpregs_28__1_), .B(
        decode_regfile_fpregs_29__1_), .S(n12961), .Z(n11952) );
  MUX2_X2 U16402 ( .A(n11952), .B(n11951), .S(n13044), .Z(n11953) );
  MUX2_X2 U16403 ( .A(decode_regfile_fpregs_26__1_), .B(
        decode_regfile_fpregs_27__1_), .S(n12961), .Z(n11954) );
  MUX2_X2 U16404 ( .A(decode_regfile_fpregs_24__1_), .B(
        decode_regfile_fpregs_25__1_), .S(n12961), .Z(n11955) );
  MUX2_X2 U16405 ( .A(n11955), .B(n11954), .S(n13044), .Z(n11956) );
  MUX2_X2 U16406 ( .A(n11956), .B(n11953), .S(n13073), .Z(n11957) );
  MUX2_X2 U16407 ( .A(decode_regfile_fpregs_22__1_), .B(
        decode_regfile_fpregs_23__1_), .S(n12961), .Z(n11958) );
  MUX2_X2 U16408 ( .A(decode_regfile_fpregs_20__1_), .B(
        decode_regfile_fpregs_21__1_), .S(n12961), .Z(n11959) );
  MUX2_X2 U16409 ( .A(n11959), .B(n11958), .S(n13044), .Z(n11960) );
  MUX2_X2 U16410 ( .A(decode_regfile_fpregs_18__1_), .B(
        decode_regfile_fpregs_19__1_), .S(n12961), .Z(n11961) );
  MUX2_X2 U16411 ( .A(decode_regfile_fpregs_16__1_), .B(
        decode_regfile_fpregs_17__1_), .S(n12961), .Z(n11962) );
  MUX2_X2 U16412 ( .A(n11962), .B(n11961), .S(n13044), .Z(n11963) );
  MUX2_X2 U16413 ( .A(n11963), .B(n11960), .S(n13073), .Z(n11964) );
  MUX2_X2 U16414 ( .A(n11964), .B(n11957), .S(n13089), .Z(n11965) );
  MUX2_X2 U16415 ( .A(decode_regfile_fpregs_14__1_), .B(
        decode_regfile_fpregs_15__1_), .S(n12961), .Z(n11966) );
  MUX2_X2 U16416 ( .A(decode_regfile_fpregs_12__1_), .B(
        decode_regfile_fpregs_13__1_), .S(n12961), .Z(n11967) );
  MUX2_X2 U16417 ( .A(n11967), .B(n11966), .S(n13044), .Z(n11968) );
  MUX2_X2 U16418 ( .A(decode_regfile_fpregs_10__1_), .B(
        decode_regfile_fpregs_11__1_), .S(n12961), .Z(n11969) );
  MUX2_X2 U16419 ( .A(decode_regfile_fpregs_8__1_), .B(
        decode_regfile_fpregs_9__1_), .S(n12961), .Z(n11970) );
  MUX2_X2 U16420 ( .A(n11970), .B(n11969), .S(n13044), .Z(n11971) );
  MUX2_X2 U16421 ( .A(n11971), .B(n11968), .S(n13073), .Z(n11972) );
  MUX2_X2 U16422 ( .A(decode_regfile_fpregs_6__1_), .B(
        decode_regfile_fpregs_7__1_), .S(n12962), .Z(n11973) );
  MUX2_X2 U16423 ( .A(decode_regfile_fpregs_4__1_), .B(
        decode_regfile_fpregs_5__1_), .S(n12962), .Z(n11974) );
  MUX2_X2 U16424 ( .A(n11974), .B(n11973), .S(n13045), .Z(n11975) );
  MUX2_X2 U16425 ( .A(decode_regfile_fpregs_2__1_), .B(
        decode_regfile_fpregs_3__1_), .S(n12962), .Z(n11976) );
  MUX2_X2 U16426 ( .A(decode_regfile_fpregs_0__1_), .B(
        decode_regfile_fpregs_1__1_), .S(n12962), .Z(n11977) );
  MUX2_X2 U16427 ( .A(n11977), .B(n11976), .S(n13045), .Z(n11978) );
  MUX2_X2 U16428 ( .A(n11978), .B(n11975), .S(n13074), .Z(n11979) );
  MUX2_X2 U16429 ( .A(n11979), .B(n11972), .S(n13089), .Z(n11980) );
  MUX2_X2 U16430 ( .A(n11980), .B(n11965), .S(n13099), .Z(decode_regfile_N162)
         );
  MUX2_X2 U16431 ( .A(decode_regfile_fpregs_30__2_), .B(
        decode_regfile_fpregs_31__2_), .S(n12962), .Z(n11981) );
  MUX2_X2 U16432 ( .A(decode_regfile_fpregs_28__2_), .B(
        decode_regfile_fpregs_29__2_), .S(n12962), .Z(n11982) );
  MUX2_X2 U16433 ( .A(n11982), .B(n11981), .S(n13045), .Z(n11983) );
  MUX2_X2 U16434 ( .A(decode_regfile_fpregs_26__2_), .B(
        decode_regfile_fpregs_27__2_), .S(n12962), .Z(n11984) );
  MUX2_X2 U16435 ( .A(decode_regfile_fpregs_24__2_), .B(
        decode_regfile_fpregs_25__2_), .S(n12962), .Z(n11985) );
  MUX2_X2 U16436 ( .A(n11985), .B(n11984), .S(n13045), .Z(n11986) );
  MUX2_X2 U16437 ( .A(n11986), .B(n11983), .S(n13074), .Z(n11987) );
  MUX2_X2 U16438 ( .A(decode_regfile_fpregs_22__2_), .B(
        decode_regfile_fpregs_23__2_), .S(n12962), .Z(n11988) );
  MUX2_X2 U16439 ( .A(decode_regfile_fpregs_20__2_), .B(
        decode_regfile_fpregs_21__2_), .S(n12962), .Z(n11989) );
  MUX2_X2 U16440 ( .A(n11989), .B(n11988), .S(n13045), .Z(n11990) );
  MUX2_X2 U16441 ( .A(decode_regfile_fpregs_18__2_), .B(
        decode_regfile_fpregs_19__2_), .S(n12962), .Z(n11991) );
  MUX2_X2 U16442 ( .A(decode_regfile_fpregs_16__2_), .B(
        decode_regfile_fpregs_17__2_), .S(n12963), .Z(n11992) );
  MUX2_X2 U16443 ( .A(n11992), .B(n11991), .S(n13045), .Z(n11993) );
  MUX2_X2 U16444 ( .A(n11993), .B(n11990), .S(n13074), .Z(n11994) );
  MUX2_X2 U16445 ( .A(n11994), .B(n11987), .S(n13089), .Z(n11995) );
  MUX2_X2 U16446 ( .A(decode_regfile_fpregs_14__2_), .B(
        decode_regfile_fpregs_15__2_), .S(n12963), .Z(n11996) );
  MUX2_X2 U16447 ( .A(decode_regfile_fpregs_12__2_), .B(
        decode_regfile_fpregs_13__2_), .S(n12963), .Z(n11997) );
  MUX2_X2 U16448 ( .A(n11997), .B(n11996), .S(n13045), .Z(n11998) );
  MUX2_X2 U16449 ( .A(decode_regfile_fpregs_10__2_), .B(
        decode_regfile_fpregs_11__2_), .S(n12963), .Z(n11999) );
  MUX2_X2 U16450 ( .A(decode_regfile_fpregs_8__2_), .B(
        decode_regfile_fpregs_9__2_), .S(n12963), .Z(n12000) );
  MUX2_X2 U16451 ( .A(n12000), .B(n11999), .S(n13045), .Z(n12001) );
  MUX2_X2 U16452 ( .A(n12001), .B(n11998), .S(n13074), .Z(n12002) );
  MUX2_X2 U16453 ( .A(decode_regfile_fpregs_6__2_), .B(
        decode_regfile_fpregs_7__2_), .S(n12963), .Z(n12003) );
  MUX2_X2 U16454 ( .A(decode_regfile_fpregs_4__2_), .B(
        decode_regfile_fpregs_5__2_), .S(n12963), .Z(n12004) );
  MUX2_X2 U16455 ( .A(n12004), .B(n12003), .S(n13045), .Z(n12005) );
  MUX2_X2 U16456 ( .A(decode_regfile_fpregs_2__2_), .B(
        decode_regfile_fpregs_3__2_), .S(n12963), .Z(n12006) );
  MUX2_X2 U16457 ( .A(decode_regfile_fpregs_0__2_), .B(
        decode_regfile_fpregs_1__2_), .S(n12963), .Z(n12007) );
  MUX2_X2 U16458 ( .A(n12007), .B(n12006), .S(n13045), .Z(n12008) );
  MUX2_X2 U16459 ( .A(n12008), .B(n12005), .S(n13074), .Z(n12009) );
  MUX2_X2 U16460 ( .A(n12009), .B(n12002), .S(n13089), .Z(n12010) );
  MUX2_X2 U16461 ( .A(n12010), .B(n11995), .S(n13099), .Z(decode_regfile_N161)
         );
  MUX2_X2 U16462 ( .A(decode_regfile_fpregs_30__3_), .B(
        decode_regfile_fpregs_31__3_), .S(n12963), .Z(n12011) );
  MUX2_X2 U16463 ( .A(decode_regfile_fpregs_28__3_), .B(
        decode_regfile_fpregs_29__3_), .S(n12963), .Z(n12012) );
  MUX2_X2 U16464 ( .A(n12012), .B(n12011), .S(n13045), .Z(n12013) );
  MUX2_X2 U16465 ( .A(decode_regfile_fpregs_26__3_), .B(
        decode_regfile_fpregs_27__3_), .S(n12964), .Z(n12014) );
  MUX2_X2 U16466 ( .A(decode_regfile_fpregs_24__3_), .B(
        decode_regfile_fpregs_25__3_), .S(n12964), .Z(n12015) );
  MUX2_X2 U16467 ( .A(n12015), .B(n12014), .S(n13046), .Z(n12016) );
  MUX2_X2 U16468 ( .A(n12016), .B(n12013), .S(n13074), .Z(n12017) );
  MUX2_X2 U16469 ( .A(decode_regfile_fpregs_22__3_), .B(
        decode_regfile_fpregs_23__3_), .S(n12964), .Z(n12018) );
  MUX2_X2 U16470 ( .A(decode_regfile_fpregs_20__3_), .B(
        decode_regfile_fpregs_21__3_), .S(n12964), .Z(n12019) );
  MUX2_X2 U16471 ( .A(n12019), .B(n12018), .S(n13046), .Z(n12020) );
  MUX2_X2 U16472 ( .A(decode_regfile_fpregs_18__3_), .B(
        decode_regfile_fpregs_19__3_), .S(n12964), .Z(n12021) );
  MUX2_X2 U16473 ( .A(decode_regfile_fpregs_16__3_), .B(
        decode_regfile_fpregs_17__3_), .S(n12964), .Z(n12022) );
  MUX2_X2 U16474 ( .A(n12022), .B(n12021), .S(n13046), .Z(n12023) );
  MUX2_X2 U16475 ( .A(n12023), .B(n12020), .S(n13074), .Z(n12024) );
  MUX2_X2 U16476 ( .A(n12024), .B(n12017), .S(n13089), .Z(n12025) );
  MUX2_X2 U16477 ( .A(decode_regfile_fpregs_14__3_), .B(
        decode_regfile_fpregs_15__3_), .S(n12964), .Z(n12026) );
  MUX2_X2 U16478 ( .A(decode_regfile_fpregs_12__3_), .B(
        decode_regfile_fpregs_13__3_), .S(n12964), .Z(n12027) );
  MUX2_X2 U16479 ( .A(n12027), .B(n12026), .S(n13046), .Z(n12028) );
  MUX2_X2 U16480 ( .A(decode_regfile_fpregs_10__3_), .B(
        decode_regfile_fpregs_11__3_), .S(n12964), .Z(n12029) );
  MUX2_X2 U16481 ( .A(decode_regfile_fpregs_8__3_), .B(
        decode_regfile_fpregs_9__3_), .S(n12964), .Z(n12030) );
  MUX2_X2 U16482 ( .A(n12030), .B(n12029), .S(n13046), .Z(n12031) );
  MUX2_X2 U16483 ( .A(n12031), .B(n12028), .S(n13074), .Z(n12032) );
  MUX2_X2 U16484 ( .A(decode_regfile_fpregs_6__3_), .B(
        decode_regfile_fpregs_7__3_), .S(n12964), .Z(n12033) );
  MUX2_X2 U16485 ( .A(decode_regfile_fpregs_4__3_), .B(
        decode_regfile_fpregs_5__3_), .S(n12965), .Z(n12034) );
  MUX2_X2 U16486 ( .A(n12034), .B(n12033), .S(n13046), .Z(n12035) );
  MUX2_X2 U16487 ( .A(decode_regfile_fpregs_2__3_), .B(
        decode_regfile_fpregs_3__3_), .S(n12965), .Z(n12036) );
  MUX2_X2 U16488 ( .A(decode_regfile_fpregs_0__3_), .B(
        decode_regfile_fpregs_1__3_), .S(n12965), .Z(n12037) );
  MUX2_X2 U16489 ( .A(n12037), .B(n12036), .S(n13046), .Z(n12038) );
  MUX2_X2 U16490 ( .A(n12038), .B(n12035), .S(n13074), .Z(n12039) );
  MUX2_X2 U16491 ( .A(n12039), .B(n12032), .S(n13089), .Z(n12040) );
  MUX2_X2 U16492 ( .A(n12040), .B(n12025), .S(n13099), .Z(decode_regfile_N160)
         );
  MUX2_X2 U16493 ( .A(decode_regfile_fpregs_30__4_), .B(
        decode_regfile_fpregs_31__4_), .S(n12965), .Z(n12041) );
  MUX2_X2 U16494 ( .A(decode_regfile_fpregs_28__4_), .B(
        decode_regfile_fpregs_29__4_), .S(n12965), .Z(n12042) );
  MUX2_X2 U16495 ( .A(n12042), .B(n12041), .S(n13046), .Z(n12043) );
  MUX2_X2 U16496 ( .A(decode_regfile_fpregs_26__4_), .B(
        decode_regfile_fpregs_27__4_), .S(n12965), .Z(n12044) );
  MUX2_X2 U16497 ( .A(decode_regfile_fpregs_24__4_), .B(
        decode_regfile_fpregs_25__4_), .S(n12965), .Z(n12045) );
  MUX2_X2 U16498 ( .A(n12045), .B(n12044), .S(n13046), .Z(n12046) );
  MUX2_X2 U16499 ( .A(n12046), .B(n12043), .S(n13074), .Z(n12047) );
  MUX2_X2 U16500 ( .A(decode_regfile_fpregs_22__4_), .B(
        decode_regfile_fpregs_23__4_), .S(n12965), .Z(n12048) );
  MUX2_X2 U16501 ( .A(decode_regfile_fpregs_20__4_), .B(
        decode_regfile_fpregs_21__4_), .S(n12965), .Z(n12049) );
  MUX2_X2 U16502 ( .A(n12049), .B(n12048), .S(n13046), .Z(n12050) );
  MUX2_X2 U16503 ( .A(decode_regfile_fpregs_18__4_), .B(
        decode_regfile_fpregs_19__4_), .S(n12965), .Z(n12051) );
  MUX2_X2 U16504 ( .A(decode_regfile_fpregs_16__4_), .B(
        decode_regfile_fpregs_17__4_), .S(n12965), .Z(n12052) );
  MUX2_X2 U16505 ( .A(n12052), .B(n12051), .S(n13046), .Z(n12053) );
  MUX2_X2 U16506 ( .A(n12053), .B(n12050), .S(n13074), .Z(n12054) );
  MUX2_X2 U16507 ( .A(n12054), .B(n12047), .S(n13089), .Z(n12055) );
  MUX2_X2 U16508 ( .A(decode_regfile_fpregs_14__4_), .B(
        decode_regfile_fpregs_15__4_), .S(n12966), .Z(n12056) );
  MUX2_X2 U16509 ( .A(decode_regfile_fpregs_12__4_), .B(
        decode_regfile_fpregs_13__4_), .S(n12966), .Z(n12057) );
  MUX2_X2 U16510 ( .A(n12057), .B(n12056), .S(n13047), .Z(n12058) );
  MUX2_X2 U16511 ( .A(decode_regfile_fpregs_10__4_), .B(
        decode_regfile_fpregs_11__4_), .S(n12966), .Z(n12059) );
  MUX2_X2 U16512 ( .A(decode_regfile_fpregs_8__4_), .B(
        decode_regfile_fpregs_9__4_), .S(n12966), .Z(n12060) );
  MUX2_X2 U16513 ( .A(n12060), .B(n12059), .S(n13047), .Z(n12061) );
  MUX2_X2 U16514 ( .A(n12061), .B(n12058), .S(n13075), .Z(n12062) );
  MUX2_X2 U16515 ( .A(decode_regfile_fpregs_6__4_), .B(
        decode_regfile_fpregs_7__4_), .S(n12966), .Z(n12063) );
  MUX2_X2 U16516 ( .A(decode_regfile_fpregs_4__4_), .B(
        decode_regfile_fpregs_5__4_), .S(n12966), .Z(n12064) );
  MUX2_X2 U16517 ( .A(n12064), .B(n12063), .S(n13047), .Z(n12065) );
  MUX2_X2 U16518 ( .A(decode_regfile_fpregs_2__4_), .B(
        decode_regfile_fpregs_3__4_), .S(n12966), .Z(n12066) );
  MUX2_X2 U16519 ( .A(decode_regfile_fpregs_0__4_), .B(
        decode_regfile_fpregs_1__4_), .S(n12966), .Z(n12067) );
  MUX2_X2 U16520 ( .A(n12067), .B(n12066), .S(n13047), .Z(n12068) );
  MUX2_X2 U16521 ( .A(n12068), .B(n12065), .S(n13075), .Z(n12069) );
  MUX2_X2 U16522 ( .A(n12069), .B(n12062), .S(n13090), .Z(n12070) );
  MUX2_X2 U16523 ( .A(n12070), .B(n12055), .S(n13099), .Z(decode_regfile_N159)
         );
  MUX2_X2 U16524 ( .A(decode_regfile_fpregs_30__5_), .B(
        decode_regfile_fpregs_31__5_), .S(n12966), .Z(n12071) );
  MUX2_X2 U16525 ( .A(decode_regfile_fpregs_28__5_), .B(
        decode_regfile_fpregs_29__5_), .S(n12966), .Z(n12072) );
  MUX2_X2 U16526 ( .A(n12072), .B(n12071), .S(n13047), .Z(n12073) );
  MUX2_X2 U16527 ( .A(decode_regfile_fpregs_26__5_), .B(
        decode_regfile_fpregs_27__5_), .S(n12966), .Z(n12074) );
  MUX2_X2 U16528 ( .A(decode_regfile_fpregs_24__5_), .B(
        decode_regfile_fpregs_25__5_), .S(n12967), .Z(n12075) );
  MUX2_X2 U16529 ( .A(n12075), .B(n12074), .S(n13047), .Z(n12076) );
  MUX2_X2 U16530 ( .A(n12076), .B(n12073), .S(n13075), .Z(n12077) );
  MUX2_X2 U16531 ( .A(decode_regfile_fpregs_22__5_), .B(
        decode_regfile_fpregs_23__5_), .S(n12967), .Z(n12078) );
  MUX2_X2 U16532 ( .A(decode_regfile_fpregs_20__5_), .B(
        decode_regfile_fpregs_21__5_), .S(n12967), .Z(n12079) );
  MUX2_X2 U16533 ( .A(n12079), .B(n12078), .S(n13047), .Z(n12080) );
  MUX2_X2 U16534 ( .A(decode_regfile_fpregs_18__5_), .B(
        decode_regfile_fpregs_19__5_), .S(n12967), .Z(n12081) );
  MUX2_X2 U16535 ( .A(decode_regfile_fpregs_16__5_), .B(
        decode_regfile_fpregs_17__5_), .S(n12967), .Z(n12082) );
  MUX2_X2 U16536 ( .A(n12082), .B(n12081), .S(n13047), .Z(n12083) );
  MUX2_X2 U16537 ( .A(n12083), .B(n12080), .S(n13075), .Z(n12084) );
  MUX2_X2 U16538 ( .A(n12084), .B(n12077), .S(n13090), .Z(n12085) );
  MUX2_X2 U16539 ( .A(decode_regfile_fpregs_14__5_), .B(
        decode_regfile_fpregs_15__5_), .S(n12967), .Z(n12086) );
  MUX2_X2 U16540 ( .A(decode_regfile_fpregs_12__5_), .B(
        decode_regfile_fpregs_13__5_), .S(n12967), .Z(n12087) );
  MUX2_X2 U16541 ( .A(n12087), .B(n12086), .S(n13047), .Z(n12088) );
  MUX2_X2 U16542 ( .A(decode_regfile_fpregs_10__5_), .B(
        decode_regfile_fpregs_11__5_), .S(n12967), .Z(n12089) );
  MUX2_X2 U16543 ( .A(decode_regfile_fpregs_8__5_), .B(
        decode_regfile_fpregs_9__5_), .S(n12967), .Z(n12090) );
  MUX2_X2 U16544 ( .A(n12090), .B(n12089), .S(n13047), .Z(n12091) );
  MUX2_X2 U16545 ( .A(n12091), .B(n12088), .S(n13075), .Z(n12092) );
  MUX2_X2 U16546 ( .A(decode_regfile_fpregs_6__5_), .B(
        decode_regfile_fpregs_7__5_), .S(n12967), .Z(n12093) );
  MUX2_X2 U16547 ( .A(decode_regfile_fpregs_4__5_), .B(
        decode_regfile_fpregs_5__5_), .S(n12967), .Z(n12094) );
  MUX2_X2 U16548 ( .A(n12094), .B(n12093), .S(n13047), .Z(n12095) );
  MUX2_X2 U16549 ( .A(decode_regfile_fpregs_2__5_), .B(
        decode_regfile_fpregs_3__5_), .S(n12968), .Z(n12096) );
  MUX2_X2 U16550 ( .A(decode_regfile_fpregs_0__5_), .B(
        decode_regfile_fpregs_1__5_), .S(n12968), .Z(n12097) );
  MUX2_X2 U16551 ( .A(n12097), .B(n12096), .S(n13048), .Z(n12098) );
  MUX2_X2 U16552 ( .A(n12098), .B(n12095), .S(n13075), .Z(n12099) );
  MUX2_X2 U16553 ( .A(n12099), .B(n12092), .S(n13090), .Z(n12100) );
  MUX2_X2 U16554 ( .A(n12100), .B(n12085), .S(n13099), .Z(decode_regfile_N158)
         );
  MUX2_X2 U16555 ( .A(decode_regfile_fpregs_30__6_), .B(
        decode_regfile_fpregs_31__6_), .S(n12968), .Z(n12101) );
  MUX2_X2 U16556 ( .A(decode_regfile_fpregs_28__6_), .B(
        decode_regfile_fpregs_29__6_), .S(n12968), .Z(n12102) );
  MUX2_X2 U16557 ( .A(n12102), .B(n12101), .S(n13048), .Z(n12103) );
  MUX2_X2 U16558 ( .A(decode_regfile_fpregs_26__6_), .B(
        decode_regfile_fpregs_27__6_), .S(n12968), .Z(n12104) );
  MUX2_X2 U16559 ( .A(decode_regfile_fpregs_24__6_), .B(
        decode_regfile_fpregs_25__6_), .S(n12968), .Z(n12105) );
  MUX2_X2 U16560 ( .A(n12105), .B(n12104), .S(n13048), .Z(n12106) );
  MUX2_X2 U16561 ( .A(n12106), .B(n12103), .S(n13075), .Z(n12107) );
  MUX2_X2 U16562 ( .A(decode_regfile_fpregs_22__6_), .B(
        decode_regfile_fpregs_23__6_), .S(n12968), .Z(n12108) );
  MUX2_X2 U16563 ( .A(decode_regfile_fpregs_20__6_), .B(
        decode_regfile_fpregs_21__6_), .S(n12968), .Z(n12109) );
  MUX2_X2 U16564 ( .A(n12109), .B(n12108), .S(n13048), .Z(n12110) );
  MUX2_X2 U16565 ( .A(decode_regfile_fpregs_18__6_), .B(
        decode_regfile_fpregs_19__6_), .S(n12968), .Z(n12111) );
  MUX2_X2 U16566 ( .A(decode_regfile_fpregs_16__6_), .B(
        decode_regfile_fpregs_17__6_), .S(n12968), .Z(n12112) );
  MUX2_X2 U16567 ( .A(n12112), .B(n12111), .S(n13048), .Z(n12113) );
  MUX2_X2 U16568 ( .A(n12113), .B(n12110), .S(n13075), .Z(n12114) );
  MUX2_X2 U16569 ( .A(n12114), .B(n12107), .S(n13090), .Z(n12115) );
  MUX2_X2 U16570 ( .A(decode_regfile_fpregs_14__6_), .B(
        decode_regfile_fpregs_15__6_), .S(n12968), .Z(n12116) );
  MUX2_X2 U16571 ( .A(decode_regfile_fpregs_12__6_), .B(
        decode_regfile_fpregs_13__6_), .S(n12969), .Z(n12117) );
  MUX2_X2 U16572 ( .A(n12117), .B(n12116), .S(n13048), .Z(n12118) );
  MUX2_X2 U16573 ( .A(decode_regfile_fpregs_10__6_), .B(
        decode_regfile_fpregs_11__6_), .S(n12969), .Z(n12119) );
  MUX2_X2 U16574 ( .A(decode_regfile_fpregs_8__6_), .B(
        decode_regfile_fpregs_9__6_), .S(n12969), .Z(n12120) );
  MUX2_X2 U16575 ( .A(n12120), .B(n12119), .S(n13048), .Z(n12121) );
  MUX2_X2 U16576 ( .A(n12121), .B(n12118), .S(n13075), .Z(n12122) );
  MUX2_X2 U16577 ( .A(decode_regfile_fpregs_6__6_), .B(
        decode_regfile_fpregs_7__6_), .S(n12969), .Z(n12123) );
  MUX2_X2 U16578 ( .A(decode_regfile_fpregs_4__6_), .B(
        decode_regfile_fpregs_5__6_), .S(n12969), .Z(n12124) );
  MUX2_X2 U16579 ( .A(n12124), .B(n12123), .S(n13048), .Z(n12125) );
  MUX2_X2 U16580 ( .A(decode_regfile_fpregs_2__6_), .B(
        decode_regfile_fpregs_3__6_), .S(n12969), .Z(n12126) );
  MUX2_X2 U16581 ( .A(decode_regfile_fpregs_0__6_), .B(
        decode_regfile_fpregs_1__6_), .S(n12969), .Z(n12127) );
  MUX2_X2 U16582 ( .A(n12127), .B(n12126), .S(n13048), .Z(n12128) );
  MUX2_X2 U16583 ( .A(n12128), .B(n12125), .S(n13075), .Z(n12129) );
  MUX2_X2 U16584 ( .A(n12129), .B(n12122), .S(n13090), .Z(n12130) );
  MUX2_X2 U16585 ( .A(n12130), .B(n12115), .S(n13099), .Z(decode_regfile_N157)
         );
  MUX2_X2 U16586 ( .A(decode_regfile_fpregs_30__7_), .B(
        decode_regfile_fpregs_31__7_), .S(n12969), .Z(n12131) );
  MUX2_X2 U16587 ( .A(decode_regfile_fpregs_28__7_), .B(
        decode_regfile_fpregs_29__7_), .S(n12969), .Z(n12132) );
  MUX2_X2 U16588 ( .A(n12132), .B(n12131), .S(n13048), .Z(n12133) );
  MUX2_X2 U16589 ( .A(decode_regfile_fpregs_26__7_), .B(
        decode_regfile_fpregs_27__7_), .S(n12969), .Z(n12134) );
  MUX2_X2 U16590 ( .A(decode_regfile_fpregs_24__7_), .B(
        decode_regfile_fpregs_25__7_), .S(n12969), .Z(n12135) );
  MUX2_X2 U16591 ( .A(n12135), .B(n12134), .S(n13048), .Z(n12136) );
  MUX2_X2 U16592 ( .A(n12136), .B(n12133), .S(n13075), .Z(n12137) );
  MUX2_X2 U16593 ( .A(decode_regfile_fpregs_22__7_), .B(
        decode_regfile_fpregs_23__7_), .S(n12970), .Z(n12138) );
  MUX2_X2 U16594 ( .A(decode_regfile_fpregs_20__7_), .B(
        decode_regfile_fpregs_21__7_), .S(n12970), .Z(n12139) );
  MUX2_X2 U16595 ( .A(n12139), .B(n12138), .S(n13049), .Z(n12140) );
  MUX2_X2 U16596 ( .A(decode_regfile_fpregs_18__7_), .B(
        decode_regfile_fpregs_19__7_), .S(n12970), .Z(n12141) );
  MUX2_X2 U16597 ( .A(decode_regfile_fpregs_16__7_), .B(
        decode_regfile_fpregs_17__7_), .S(n12970), .Z(n12142) );
  MUX2_X2 U16598 ( .A(n12142), .B(n12141), .S(n13049), .Z(n12143) );
  MUX2_X2 U16599 ( .A(n12143), .B(n12140), .S(n13076), .Z(n12144) );
  MUX2_X2 U16600 ( .A(n12144), .B(n12137), .S(n13090), .Z(n12145) );
  MUX2_X2 U16601 ( .A(decode_regfile_fpregs_14__7_), .B(
        decode_regfile_fpregs_15__7_), .S(n12970), .Z(n12146) );
  MUX2_X2 U16602 ( .A(decode_regfile_fpregs_12__7_), .B(
        decode_regfile_fpregs_13__7_), .S(n12970), .Z(n12147) );
  MUX2_X2 U16603 ( .A(n12147), .B(n12146), .S(n13049), .Z(n12148) );
  MUX2_X2 U16604 ( .A(decode_regfile_fpregs_10__7_), .B(
        decode_regfile_fpregs_11__7_), .S(n12970), .Z(n12149) );
  MUX2_X2 U16605 ( .A(decode_regfile_fpregs_8__7_), .B(
        decode_regfile_fpregs_9__7_), .S(n12970), .Z(n12150) );
  MUX2_X2 U16606 ( .A(n12150), .B(n12149), .S(n13049), .Z(n12151) );
  MUX2_X2 U16607 ( .A(n12151), .B(n12148), .S(n13076), .Z(n12152) );
  MUX2_X2 U16608 ( .A(decode_regfile_fpregs_6__7_), .B(
        decode_regfile_fpregs_7__7_), .S(n12970), .Z(n12153) );
  MUX2_X2 U16609 ( .A(decode_regfile_fpregs_4__7_), .B(
        decode_regfile_fpregs_5__7_), .S(n12970), .Z(n12154) );
  MUX2_X2 U16610 ( .A(n12154), .B(n12153), .S(n13049), .Z(n12155) );
  MUX2_X2 U16611 ( .A(decode_regfile_fpregs_2__7_), .B(
        decode_regfile_fpregs_3__7_), .S(n12970), .Z(n12156) );
  MUX2_X2 U16612 ( .A(decode_regfile_fpregs_0__7_), .B(
        decode_regfile_fpregs_1__7_), .S(n12971), .Z(n12157) );
  MUX2_X2 U16613 ( .A(n12157), .B(n12156), .S(n13049), .Z(n12158) );
  MUX2_X2 U16614 ( .A(n12158), .B(n12155), .S(n13076), .Z(n12159) );
  MUX2_X2 U16615 ( .A(n12159), .B(n12152), .S(n13090), .Z(n12160) );
  MUX2_X2 U16616 ( .A(n12160), .B(n12145), .S(n13099), .Z(decode_regfile_N156)
         );
  MUX2_X2 U16617 ( .A(decode_regfile_fpregs_30__8_), .B(
        decode_regfile_fpregs_31__8_), .S(n12971), .Z(n12161) );
  MUX2_X2 U16618 ( .A(decode_regfile_fpregs_28__8_), .B(
        decode_regfile_fpregs_29__8_), .S(n12971), .Z(n12162) );
  MUX2_X2 U16619 ( .A(n12162), .B(n12161), .S(n13049), .Z(n12163) );
  MUX2_X2 U16620 ( .A(decode_regfile_fpregs_26__8_), .B(
        decode_regfile_fpregs_27__8_), .S(n12971), .Z(n12164) );
  MUX2_X2 U16621 ( .A(decode_regfile_fpregs_24__8_), .B(
        decode_regfile_fpregs_25__8_), .S(n12971), .Z(n12165) );
  MUX2_X2 U16622 ( .A(n12165), .B(n12164), .S(n13049), .Z(n12166) );
  MUX2_X2 U16623 ( .A(n12166), .B(n12163), .S(n13076), .Z(n12167) );
  MUX2_X2 U16624 ( .A(decode_regfile_fpregs_22__8_), .B(
        decode_regfile_fpregs_23__8_), .S(n12971), .Z(n12168) );
  MUX2_X2 U16625 ( .A(decode_regfile_fpregs_20__8_), .B(
        decode_regfile_fpregs_21__8_), .S(n12971), .Z(n12169) );
  MUX2_X2 U16626 ( .A(n12169), .B(n12168), .S(n13049), .Z(n12170) );
  MUX2_X2 U16627 ( .A(decode_regfile_fpregs_18__8_), .B(
        decode_regfile_fpregs_19__8_), .S(n12971), .Z(n12171) );
  MUX2_X2 U16628 ( .A(decode_regfile_fpregs_16__8_), .B(
        decode_regfile_fpregs_17__8_), .S(n12971), .Z(n12172) );
  MUX2_X2 U16629 ( .A(n12172), .B(n12171), .S(n13049), .Z(n12173) );
  MUX2_X2 U16630 ( .A(n12173), .B(n12170), .S(n13076), .Z(n12174) );
  MUX2_X2 U16631 ( .A(n12174), .B(n12167), .S(n13090), .Z(n12175) );
  MUX2_X2 U16632 ( .A(decode_regfile_fpregs_14__8_), .B(
        decode_regfile_fpregs_15__8_), .S(n12971), .Z(n12176) );
  MUX2_X2 U16633 ( .A(decode_regfile_fpregs_12__8_), .B(
        decode_regfile_fpregs_13__8_), .S(n12971), .Z(n12177) );
  MUX2_X2 U16634 ( .A(n12177), .B(n12176), .S(n13049), .Z(n12178) );
  MUX2_X2 U16635 ( .A(decode_regfile_fpregs_10__8_), .B(
        decode_regfile_fpregs_11__8_), .S(n12972), .Z(n12179) );
  MUX2_X2 U16636 ( .A(decode_regfile_fpregs_8__8_), .B(
        decode_regfile_fpregs_9__8_), .S(n12972), .Z(n12180) );
  MUX2_X2 U16637 ( .A(n12180), .B(n12179), .S(n13050), .Z(n12181) );
  MUX2_X2 U16638 ( .A(n12181), .B(n12178), .S(n13076), .Z(n12182) );
  MUX2_X2 U16639 ( .A(decode_regfile_fpregs_6__8_), .B(
        decode_regfile_fpregs_7__8_), .S(n12972), .Z(n12183) );
  MUX2_X2 U16640 ( .A(decode_regfile_fpregs_4__8_), .B(
        decode_regfile_fpregs_5__8_), .S(n12972), .Z(n12184) );
  MUX2_X2 U16641 ( .A(n12184), .B(n12183), .S(n13050), .Z(n12185) );
  MUX2_X2 U16642 ( .A(decode_regfile_fpregs_2__8_), .B(
        decode_regfile_fpregs_3__8_), .S(n12972), .Z(n12186) );
  MUX2_X2 U16643 ( .A(decode_regfile_fpregs_0__8_), .B(
        decode_regfile_fpregs_1__8_), .S(n12972), .Z(n12187) );
  MUX2_X2 U16644 ( .A(n12187), .B(n12186), .S(n13050), .Z(n12188) );
  MUX2_X2 U16645 ( .A(n12188), .B(n12185), .S(n13076), .Z(n12189) );
  MUX2_X2 U16646 ( .A(n12189), .B(n12182), .S(n13090), .Z(n12190) );
  MUX2_X2 U16647 ( .A(n12190), .B(n12175), .S(n13099), .Z(decode_regfile_N155)
         );
  MUX2_X2 U16648 ( .A(decode_regfile_fpregs_30__9_), .B(
        decode_regfile_fpregs_31__9_), .S(n12972), .Z(n12191) );
  MUX2_X2 U16649 ( .A(decode_regfile_fpregs_28__9_), .B(
        decode_regfile_fpregs_29__9_), .S(n12972), .Z(n12192) );
  MUX2_X2 U16650 ( .A(n12192), .B(n12191), .S(n13050), .Z(n12193) );
  MUX2_X2 U16651 ( .A(decode_regfile_fpregs_26__9_), .B(
        decode_regfile_fpregs_27__9_), .S(n12972), .Z(n12194) );
  MUX2_X2 U16652 ( .A(decode_regfile_fpregs_24__9_), .B(
        decode_regfile_fpregs_25__9_), .S(n12972), .Z(n12195) );
  MUX2_X2 U16653 ( .A(n12195), .B(n12194), .S(n13050), .Z(n12196) );
  MUX2_X2 U16654 ( .A(n12196), .B(n12193), .S(n13076), .Z(n12197) );
  MUX2_X2 U16655 ( .A(decode_regfile_fpregs_22__9_), .B(
        decode_regfile_fpregs_23__9_), .S(n12972), .Z(n12198) );
  MUX2_X2 U16656 ( .A(decode_regfile_fpregs_20__9_), .B(
        decode_regfile_fpregs_21__9_), .S(n12973), .Z(n12199) );
  MUX2_X2 U16657 ( .A(n12199), .B(n12198), .S(n13050), .Z(n12200) );
  MUX2_X2 U16658 ( .A(decode_regfile_fpregs_18__9_), .B(
        decode_regfile_fpregs_19__9_), .S(n12973), .Z(n12201) );
  MUX2_X2 U16659 ( .A(decode_regfile_fpregs_16__9_), .B(
        decode_regfile_fpregs_17__9_), .S(n12973), .Z(n12202) );
  MUX2_X2 U16660 ( .A(n12202), .B(n12201), .S(n13050), .Z(n12203) );
  MUX2_X2 U16661 ( .A(n12203), .B(n12200), .S(n13076), .Z(n12204) );
  MUX2_X2 U16662 ( .A(n12204), .B(n12197), .S(n13090), .Z(n12205) );
  MUX2_X2 U16663 ( .A(decode_regfile_fpregs_14__9_), .B(
        decode_regfile_fpregs_15__9_), .S(n12973), .Z(n12206) );
  MUX2_X2 U16664 ( .A(decode_regfile_fpregs_12__9_), .B(
        decode_regfile_fpregs_13__9_), .S(n12973), .Z(n12207) );
  MUX2_X2 U16665 ( .A(n12207), .B(n12206), .S(n13050), .Z(n12208) );
  MUX2_X2 U16666 ( .A(decode_regfile_fpregs_10__9_), .B(
        decode_regfile_fpregs_11__9_), .S(n12973), .Z(n12209) );
  MUX2_X2 U16667 ( .A(decode_regfile_fpregs_8__9_), .B(
        decode_regfile_fpregs_9__9_), .S(n12973), .Z(n12210) );
  MUX2_X2 U16668 ( .A(n12210), .B(n12209), .S(n13050), .Z(n12211) );
  MUX2_X2 U16669 ( .A(n12211), .B(n12208), .S(n13076), .Z(n12212) );
  MUX2_X2 U16670 ( .A(decode_regfile_fpregs_6__9_), .B(
        decode_regfile_fpregs_7__9_), .S(n12973), .Z(n12213) );
  MUX2_X2 U16671 ( .A(decode_regfile_fpregs_4__9_), .B(
        decode_regfile_fpregs_5__9_), .S(n12973), .Z(n12214) );
  MUX2_X2 U16672 ( .A(n12214), .B(n12213), .S(n13050), .Z(n12215) );
  MUX2_X2 U16673 ( .A(decode_regfile_fpregs_2__9_), .B(
        decode_regfile_fpregs_3__9_), .S(n12973), .Z(n12216) );
  MUX2_X2 U16674 ( .A(decode_regfile_fpregs_0__9_), .B(
        decode_regfile_fpregs_1__9_), .S(n12973), .Z(n12217) );
  MUX2_X2 U16675 ( .A(n12217), .B(n12216), .S(n13050), .Z(n12218) );
  MUX2_X2 U16676 ( .A(n12218), .B(n12215), .S(n13076), .Z(n12219) );
  MUX2_X2 U16677 ( .A(n12219), .B(n12212), .S(n13090), .Z(n12220) );
  MUX2_X2 U16678 ( .A(n12220), .B(n12205), .S(n13099), .Z(decode_regfile_N154)
         );
  MUX2_X2 U16679 ( .A(decode_regfile_fpregs_30__10_), .B(
        decode_regfile_fpregs_31__10_), .S(n12974), .Z(n12221) );
  MUX2_X2 U16680 ( .A(decode_regfile_fpregs_28__10_), .B(
        decode_regfile_fpregs_29__10_), .S(n12974), .Z(n12222) );
  MUX2_X2 U16681 ( .A(n12222), .B(n12221), .S(n13051), .Z(n12223) );
  MUX2_X2 U16682 ( .A(decode_regfile_fpregs_26__10_), .B(
        decode_regfile_fpregs_27__10_), .S(n12974), .Z(n12224) );
  MUX2_X2 U16683 ( .A(decode_regfile_fpregs_24__10_), .B(
        decode_regfile_fpregs_25__10_), .S(n12974), .Z(n12225) );
  MUX2_X2 U16684 ( .A(n12225), .B(n12224), .S(n13051), .Z(n12226) );
  MUX2_X2 U16685 ( .A(n12226), .B(n12223), .S(n13077), .Z(n12227) );
  MUX2_X2 U16686 ( .A(decode_regfile_fpregs_22__10_), .B(
        decode_regfile_fpregs_23__10_), .S(n12974), .Z(n12228) );
  MUX2_X2 U16687 ( .A(decode_regfile_fpregs_20__10_), .B(
        decode_regfile_fpregs_21__10_), .S(n12974), .Z(n12229) );
  MUX2_X2 U16688 ( .A(n12229), .B(n12228), .S(n13051), .Z(n12230) );
  MUX2_X2 U16689 ( .A(decode_regfile_fpregs_18__10_), .B(
        decode_regfile_fpregs_19__10_), .S(n12974), .Z(n12231) );
  MUX2_X2 U16690 ( .A(decode_regfile_fpregs_16__10_), .B(
        decode_regfile_fpregs_17__10_), .S(n12974), .Z(n12232) );
  MUX2_X2 U16691 ( .A(n12232), .B(n12231), .S(n13051), .Z(n12233) );
  MUX2_X2 U16692 ( .A(n12233), .B(n12230), .S(n13077), .Z(n12234) );
  MUX2_X2 U16693 ( .A(n12234), .B(n12227), .S(n13091), .Z(n12235) );
  MUX2_X2 U16694 ( .A(decode_regfile_fpregs_14__10_), .B(
        decode_regfile_fpregs_15__10_), .S(n12974), .Z(n12236) );
  MUX2_X2 U16695 ( .A(decode_regfile_fpregs_12__10_), .B(
        decode_regfile_fpregs_13__10_), .S(n12974), .Z(n12237) );
  MUX2_X2 U16696 ( .A(n12237), .B(n12236), .S(n13051), .Z(n12238) );
  MUX2_X2 U16697 ( .A(decode_regfile_fpregs_10__10_), .B(
        decode_regfile_fpregs_11__10_), .S(n12974), .Z(n12239) );
  MUX2_X2 U16698 ( .A(decode_regfile_fpregs_8__10_), .B(
        decode_regfile_fpregs_9__10_), .S(n12975), .Z(n12240) );
  MUX2_X2 U16699 ( .A(n12240), .B(n12239), .S(n13051), .Z(n12241) );
  MUX2_X2 U16700 ( .A(n12241), .B(n12238), .S(n13077), .Z(n12242) );
  MUX2_X2 U16701 ( .A(decode_regfile_fpregs_6__10_), .B(
        decode_regfile_fpregs_7__10_), .S(n12975), .Z(n12243) );
  MUX2_X2 U16702 ( .A(decode_regfile_fpregs_4__10_), .B(
        decode_regfile_fpregs_5__10_), .S(n12975), .Z(n12244) );
  MUX2_X2 U16703 ( .A(n12244), .B(n12243), .S(n13051), .Z(n12245) );
  MUX2_X2 U16704 ( .A(decode_regfile_fpregs_2__10_), .B(
        decode_regfile_fpregs_3__10_), .S(n12975), .Z(n12246) );
  MUX2_X2 U16705 ( .A(decode_regfile_fpregs_0__10_), .B(
        decode_regfile_fpregs_1__10_), .S(n12975), .Z(n12247) );
  MUX2_X2 U16706 ( .A(n12247), .B(n12246), .S(n13051), .Z(n12248) );
  MUX2_X2 U16707 ( .A(n12248), .B(n12245), .S(n13077), .Z(n12249) );
  MUX2_X2 U16708 ( .A(n12249), .B(n12242), .S(n13091), .Z(n12250) );
  MUX2_X2 U16709 ( .A(n12250), .B(n12235), .S(n13100), .Z(decode_regfile_N153)
         );
  MUX2_X2 U16710 ( .A(decode_regfile_fpregs_30__11_), .B(
        decode_regfile_fpregs_31__11_), .S(n12975), .Z(n12251) );
  MUX2_X2 U16711 ( .A(decode_regfile_fpregs_28__11_), .B(
        decode_regfile_fpregs_29__11_), .S(n12975), .Z(n12252) );
  MUX2_X2 U16712 ( .A(n12252), .B(n12251), .S(n13051), .Z(n12253) );
  MUX2_X2 U16713 ( .A(decode_regfile_fpregs_26__11_), .B(
        decode_regfile_fpregs_27__11_), .S(n12975), .Z(n12254) );
  MUX2_X2 U16714 ( .A(decode_regfile_fpregs_24__11_), .B(
        decode_regfile_fpregs_25__11_), .S(n12975), .Z(n12255) );
  MUX2_X2 U16715 ( .A(n12255), .B(n12254), .S(n13051), .Z(n12256) );
  MUX2_X2 U16716 ( .A(n12256), .B(n12253), .S(n13077), .Z(n12257) );
  MUX2_X2 U16717 ( .A(decode_regfile_fpregs_22__11_), .B(
        decode_regfile_fpregs_23__11_), .S(n12975), .Z(n12258) );
  MUX2_X2 U16718 ( .A(decode_regfile_fpregs_20__11_), .B(
        decode_regfile_fpregs_21__11_), .S(n12975), .Z(n12259) );
  MUX2_X2 U16719 ( .A(n12259), .B(n12258), .S(n13051), .Z(n12260) );
  MUX2_X2 U16720 ( .A(decode_regfile_fpregs_18__11_), .B(
        decode_regfile_fpregs_19__11_), .S(n12976), .Z(n12261) );
  MUX2_X2 U16721 ( .A(decode_regfile_fpregs_16__11_), .B(
        decode_regfile_fpregs_17__11_), .S(n12976), .Z(n12262) );
  MUX2_X2 U16722 ( .A(n12262), .B(n12261), .S(n13008), .Z(n12263) );
  MUX2_X2 U16723 ( .A(n12263), .B(n12260), .S(n13077), .Z(n12264) );
  MUX2_X2 U16724 ( .A(n12264), .B(n12257), .S(n13091), .Z(n12265) );
  MUX2_X2 U16725 ( .A(decode_regfile_fpregs_14__11_), .B(
        decode_regfile_fpregs_15__11_), .S(n12976), .Z(n12266) );
  MUX2_X2 U16726 ( .A(decode_regfile_fpregs_12__11_), .B(
        decode_regfile_fpregs_13__11_), .S(n12976), .Z(n12267) );
  MUX2_X2 U16727 ( .A(n12267), .B(n12266), .S(n13006), .Z(n12268) );
  MUX2_X2 U16728 ( .A(decode_regfile_fpregs_10__11_), .B(
        decode_regfile_fpregs_11__11_), .S(n12976), .Z(n12269) );
  MUX2_X2 U16729 ( .A(decode_regfile_fpregs_8__11_), .B(
        decode_regfile_fpregs_9__11_), .S(n12976), .Z(n12270) );
  MUX2_X2 U16730 ( .A(n12270), .B(n12269), .S(n13007), .Z(n12271) );
  MUX2_X2 U16731 ( .A(n12271), .B(n12268), .S(n13077), .Z(n12272) );
  MUX2_X2 U16732 ( .A(decode_regfile_fpregs_6__11_), .B(
        decode_regfile_fpregs_7__11_), .S(n12976), .Z(n12273) );
  MUX2_X2 U16733 ( .A(decode_regfile_fpregs_4__11_), .B(
        decode_regfile_fpregs_5__11_), .S(n12976), .Z(n12274) );
  MUX2_X2 U16734 ( .A(n12274), .B(n12273), .S(n13013), .Z(n12275) );
  MUX2_X2 U16735 ( .A(decode_regfile_fpregs_2__11_), .B(
        decode_regfile_fpregs_3__11_), .S(n12976), .Z(n12276) );
  MUX2_X2 U16736 ( .A(decode_regfile_fpregs_0__11_), .B(
        decode_regfile_fpregs_1__11_), .S(n12976), .Z(n12277) );
  MUX2_X2 U16737 ( .A(n12277), .B(n12276), .S(n13016), .Z(n12278) );
  MUX2_X2 U16738 ( .A(n12278), .B(n12275), .S(n13077), .Z(n12279) );
  MUX2_X2 U16739 ( .A(n12279), .B(n12272), .S(n13091), .Z(n12280) );
  MUX2_X2 U16740 ( .A(n12280), .B(n12265), .S(n13100), .Z(decode_regfile_N152)
         );
  MUX2_X2 U16741 ( .A(decode_regfile_fpregs_30__12_), .B(
        decode_regfile_fpregs_31__12_), .S(n12976), .Z(n12281) );
  MUX2_X2 U16742 ( .A(decode_regfile_fpregs_28__12_), .B(
        decode_regfile_fpregs_29__12_), .S(n12977), .Z(n12282) );
  MUX2_X2 U16743 ( .A(n12282), .B(n12281), .S(n13010), .Z(n12283) );
  MUX2_X2 U16744 ( .A(decode_regfile_fpregs_26__12_), .B(
        decode_regfile_fpregs_27__12_), .S(n12977), .Z(n12284) );
  MUX2_X2 U16745 ( .A(decode_regfile_fpregs_24__12_), .B(
        decode_regfile_fpregs_25__12_), .S(n12977), .Z(n12285) );
  MUX2_X2 U16746 ( .A(n12285), .B(n12284), .S(n13012), .Z(n12286) );
  MUX2_X2 U16747 ( .A(n12286), .B(n12283), .S(n13077), .Z(n12287) );
  MUX2_X2 U16748 ( .A(decode_regfile_fpregs_22__12_), .B(
        decode_regfile_fpregs_23__12_), .S(n12977), .Z(n12288) );
  MUX2_X2 U16749 ( .A(decode_regfile_fpregs_20__12_), .B(
        decode_regfile_fpregs_21__12_), .S(n12977), .Z(n12289) );
  MUX2_X2 U16750 ( .A(n12289), .B(n12288), .S(n13011), .Z(n12290) );
  MUX2_X2 U16751 ( .A(decode_regfile_fpregs_18__12_), .B(
        decode_regfile_fpregs_19__12_), .S(n12977), .Z(n12291) );
  MUX2_X2 U16752 ( .A(decode_regfile_fpregs_16__12_), .B(
        decode_regfile_fpregs_17__12_), .S(n12977), .Z(n12292) );
  MUX2_X2 U16753 ( .A(n12292), .B(n12291), .S(n13014), .Z(n12293) );
  MUX2_X2 U16754 ( .A(n12293), .B(n12290), .S(n13077), .Z(n12294) );
  MUX2_X2 U16755 ( .A(n12294), .B(n12287), .S(n13091), .Z(n12295) );
  MUX2_X2 U16756 ( .A(decode_regfile_fpregs_14__12_), .B(
        decode_regfile_fpregs_15__12_), .S(n12977), .Z(n12296) );
  MUX2_X2 U16757 ( .A(decode_regfile_fpregs_12__12_), .B(
        decode_regfile_fpregs_13__12_), .S(n12977), .Z(n12297) );
  MUX2_X2 U16758 ( .A(n12297), .B(n12296), .S(n13010), .Z(n12298) );
  MUX2_X2 U16759 ( .A(decode_regfile_fpregs_10__12_), .B(
        decode_regfile_fpregs_11__12_), .S(n12977), .Z(n12299) );
  MUX2_X2 U16760 ( .A(decode_regfile_fpregs_8__12_), .B(
        decode_regfile_fpregs_9__12_), .S(n12977), .Z(n12300) );
  MUX2_X2 U16761 ( .A(n12300), .B(n12299), .S(n13020), .Z(n12301) );
  MUX2_X2 U16762 ( .A(n12301), .B(n12298), .S(n13077), .Z(n12302) );
  MUX2_X2 U16763 ( .A(decode_regfile_fpregs_6__12_), .B(
        decode_regfile_fpregs_7__12_), .S(n12978), .Z(n12303) );
  MUX2_X2 U16764 ( .A(decode_regfile_fpregs_4__12_), .B(
        decode_regfile_fpregs_5__12_), .S(n12978), .Z(n12304) );
  MUX2_X2 U16765 ( .A(n12304), .B(n12303), .S(n13052), .Z(n12305) );
  MUX2_X2 U16766 ( .A(decode_regfile_fpregs_2__12_), .B(
        decode_regfile_fpregs_3__12_), .S(n12978), .Z(n12306) );
  MUX2_X2 U16767 ( .A(decode_regfile_fpregs_0__12_), .B(
        decode_regfile_fpregs_1__12_), .S(n12978), .Z(n12307) );
  MUX2_X2 U16768 ( .A(n12307), .B(n12306), .S(n13052), .Z(n12308) );
  MUX2_X2 U16769 ( .A(n12308), .B(n12305), .S(n13078), .Z(n12309) );
  MUX2_X2 U16770 ( .A(n12309), .B(n12302), .S(n13091), .Z(n12310) );
  MUX2_X2 U16771 ( .A(n12310), .B(n12295), .S(n13100), .Z(decode_regfile_N151)
         );
  MUX2_X2 U16772 ( .A(decode_regfile_fpregs_30__13_), .B(
        decode_regfile_fpregs_31__13_), .S(n12978), .Z(n12311) );
  MUX2_X2 U16773 ( .A(decode_regfile_fpregs_28__13_), .B(
        decode_regfile_fpregs_29__13_), .S(n12978), .Z(n12312) );
  MUX2_X2 U16774 ( .A(n12312), .B(n12311), .S(n13052), .Z(n12313) );
  MUX2_X2 U16775 ( .A(decode_regfile_fpregs_26__13_), .B(
        decode_regfile_fpregs_27__13_), .S(n12978), .Z(n12314) );
  MUX2_X2 U16776 ( .A(decode_regfile_fpregs_24__13_), .B(
        decode_regfile_fpregs_25__13_), .S(n12978), .Z(n12315) );
  MUX2_X2 U16777 ( .A(n12315), .B(n12314), .S(n13052), .Z(n12316) );
  MUX2_X2 U16778 ( .A(n12316), .B(n12313), .S(n13078), .Z(n12317) );
  MUX2_X2 U16779 ( .A(decode_regfile_fpregs_22__13_), .B(
        decode_regfile_fpregs_23__13_), .S(n12978), .Z(n12318) );
  MUX2_X2 U16780 ( .A(decode_regfile_fpregs_20__13_), .B(
        decode_regfile_fpregs_21__13_), .S(n12978), .Z(n12319) );
  MUX2_X2 U16781 ( .A(n12319), .B(n12318), .S(n13052), .Z(n12320) );
  MUX2_X2 U16782 ( .A(decode_regfile_fpregs_18__13_), .B(
        decode_regfile_fpregs_19__13_), .S(n12978), .Z(n12321) );
  MUX2_X2 U16783 ( .A(decode_regfile_fpregs_16__13_), .B(
        decode_regfile_fpregs_17__13_), .S(n12979), .Z(n12322) );
  MUX2_X2 U16784 ( .A(n12322), .B(n12321), .S(n13052), .Z(n12323) );
  MUX2_X2 U16785 ( .A(n12323), .B(n12320), .S(n13078), .Z(n12324) );
  MUX2_X2 U16786 ( .A(n12324), .B(n12317), .S(n13091), .Z(n12325) );
  MUX2_X2 U16787 ( .A(decode_regfile_fpregs_14__13_), .B(
        decode_regfile_fpregs_15__13_), .S(n12979), .Z(n12326) );
  MUX2_X2 U16788 ( .A(decode_regfile_fpregs_12__13_), .B(
        decode_regfile_fpregs_13__13_), .S(n12979), .Z(n12327) );
  MUX2_X2 U16789 ( .A(n12327), .B(n12326), .S(n13052), .Z(n12328) );
  MUX2_X2 U16790 ( .A(decode_regfile_fpregs_10__13_), .B(
        decode_regfile_fpregs_11__13_), .S(n12979), .Z(n12329) );
  MUX2_X2 U16791 ( .A(decode_regfile_fpregs_8__13_), .B(
        decode_regfile_fpregs_9__13_), .S(n12979), .Z(n12330) );
  MUX2_X2 U16792 ( .A(n12330), .B(n12329), .S(n13052), .Z(n12331) );
  MUX2_X2 U16793 ( .A(n12331), .B(n12328), .S(n13078), .Z(n12332) );
  MUX2_X2 U16794 ( .A(decode_regfile_fpregs_6__13_), .B(
        decode_regfile_fpregs_7__13_), .S(n12979), .Z(n12333) );
  MUX2_X2 U16795 ( .A(decode_regfile_fpregs_4__13_), .B(
        decode_regfile_fpregs_5__13_), .S(n12979), .Z(n12334) );
  MUX2_X2 U16796 ( .A(n12334), .B(n12333), .S(n13052), .Z(n12335) );
  MUX2_X2 U16797 ( .A(decode_regfile_fpregs_2__13_), .B(
        decode_regfile_fpregs_3__13_), .S(n12979), .Z(n12336) );
  MUX2_X2 U16798 ( .A(decode_regfile_fpregs_0__13_), .B(
        decode_regfile_fpregs_1__13_), .S(n12979), .Z(n12337) );
  MUX2_X2 U16799 ( .A(n12337), .B(n12336), .S(n13052), .Z(n12338) );
  MUX2_X2 U16800 ( .A(n12338), .B(n12335), .S(n13078), .Z(n12339) );
  MUX2_X2 U16801 ( .A(n12339), .B(n12332), .S(n13091), .Z(n12340) );
  MUX2_X2 U16802 ( .A(n12340), .B(n12325), .S(n13100), .Z(decode_regfile_N150)
         );
  MUX2_X2 U16803 ( .A(decode_regfile_fpregs_30__14_), .B(
        decode_regfile_fpregs_31__14_), .S(n12979), .Z(n12341) );
  MUX2_X2 U16804 ( .A(decode_regfile_fpregs_28__14_), .B(
        decode_regfile_fpregs_29__14_), .S(n12979), .Z(n12342) );
  MUX2_X2 U16805 ( .A(n12342), .B(n12341), .S(n13052), .Z(n12343) );
  MUX2_X2 U16806 ( .A(decode_regfile_fpregs_26__14_), .B(
        decode_regfile_fpregs_27__14_), .S(n12980), .Z(n12344) );
  MUX2_X2 U16807 ( .A(decode_regfile_fpregs_24__14_), .B(
        decode_regfile_fpregs_25__14_), .S(n12980), .Z(n12345) );
  MUX2_X2 U16808 ( .A(n12345), .B(n12344), .S(n13053), .Z(n12346) );
  MUX2_X2 U16809 ( .A(n12346), .B(n12343), .S(n13078), .Z(n12347) );
  MUX2_X2 U16810 ( .A(decode_regfile_fpregs_22__14_), .B(
        decode_regfile_fpregs_23__14_), .S(n12980), .Z(n12348) );
  MUX2_X2 U16811 ( .A(decode_regfile_fpregs_20__14_), .B(
        decode_regfile_fpregs_21__14_), .S(n12980), .Z(n12349) );
  MUX2_X2 U16812 ( .A(n12349), .B(n12348), .S(n13053), .Z(n12350) );
  MUX2_X2 U16813 ( .A(decode_regfile_fpregs_18__14_), .B(
        decode_regfile_fpregs_19__14_), .S(n12980), .Z(n12351) );
  MUX2_X2 U16814 ( .A(decode_regfile_fpregs_16__14_), .B(
        decode_regfile_fpregs_17__14_), .S(n12980), .Z(n12352) );
  MUX2_X2 U16815 ( .A(n12352), .B(n12351), .S(n13053), .Z(n12353) );
  MUX2_X2 U16816 ( .A(n12353), .B(n12350), .S(n13078), .Z(n12354) );
  MUX2_X2 U16817 ( .A(n12354), .B(n12347), .S(n13091), .Z(n12355) );
  MUX2_X2 U16818 ( .A(decode_regfile_fpregs_14__14_), .B(
        decode_regfile_fpregs_15__14_), .S(n12980), .Z(n12356) );
  MUX2_X2 U16819 ( .A(decode_regfile_fpregs_12__14_), .B(
        decode_regfile_fpregs_13__14_), .S(n12980), .Z(n12357) );
  MUX2_X2 U16820 ( .A(n12357), .B(n12356), .S(n13053), .Z(n12358) );
  MUX2_X2 U16821 ( .A(decode_regfile_fpregs_10__14_), .B(
        decode_regfile_fpregs_11__14_), .S(n12980), .Z(n12359) );
  MUX2_X2 U16822 ( .A(decode_regfile_fpregs_8__14_), .B(
        decode_regfile_fpregs_9__14_), .S(n12980), .Z(n12360) );
  MUX2_X2 U16823 ( .A(n12360), .B(n12359), .S(n13053), .Z(n12361) );
  MUX2_X2 U16824 ( .A(n12361), .B(n12358), .S(n13078), .Z(n12362) );
  MUX2_X2 U16825 ( .A(decode_regfile_fpregs_6__14_), .B(
        decode_regfile_fpregs_7__14_), .S(n12980), .Z(n12363) );
  MUX2_X2 U16826 ( .A(decode_regfile_fpregs_4__14_), .B(
        decode_regfile_fpregs_5__14_), .S(n12981), .Z(n12364) );
  MUX2_X2 U16827 ( .A(n12364), .B(n12363), .S(n13053), .Z(n12365) );
  MUX2_X2 U16828 ( .A(decode_regfile_fpregs_2__14_), .B(
        decode_regfile_fpregs_3__14_), .S(n12981), .Z(n12366) );
  MUX2_X2 U16829 ( .A(decode_regfile_fpregs_0__14_), .B(
        decode_regfile_fpregs_1__14_), .S(n12981), .Z(n12367) );
  MUX2_X2 U16830 ( .A(n12367), .B(n12366), .S(n13053), .Z(n12368) );
  MUX2_X2 U16831 ( .A(n12368), .B(n12365), .S(n13078), .Z(n12369) );
  MUX2_X2 U16832 ( .A(n12369), .B(n12362), .S(n13091), .Z(n12370) );
  MUX2_X2 U16833 ( .A(n12370), .B(n12355), .S(n13100), .Z(decode_regfile_N149)
         );
  MUX2_X2 U16834 ( .A(decode_regfile_fpregs_30__15_), .B(
        decode_regfile_fpregs_31__15_), .S(n12981), .Z(n12371) );
  MUX2_X2 U16835 ( .A(decode_regfile_fpregs_28__15_), .B(
        decode_regfile_fpregs_29__15_), .S(n12981), .Z(n12372) );
  MUX2_X2 U16836 ( .A(n12372), .B(n12371), .S(n13053), .Z(n12373) );
  MUX2_X2 U16837 ( .A(decode_regfile_fpregs_26__15_), .B(
        decode_regfile_fpregs_27__15_), .S(n12981), .Z(n12374) );
  MUX2_X2 U16838 ( .A(decode_regfile_fpregs_24__15_), .B(
        decode_regfile_fpregs_25__15_), .S(n12981), .Z(n12375) );
  MUX2_X2 U16839 ( .A(n12375), .B(n12374), .S(n13053), .Z(n12376) );
  MUX2_X2 U16840 ( .A(n12376), .B(n12373), .S(n13078), .Z(n12377) );
  MUX2_X2 U16841 ( .A(decode_regfile_fpregs_22__15_), .B(
        decode_regfile_fpregs_23__15_), .S(n12981), .Z(n12378) );
  MUX2_X2 U16842 ( .A(decode_regfile_fpregs_20__15_), .B(
        decode_regfile_fpregs_21__15_), .S(n12981), .Z(n12379) );
  MUX2_X2 U16843 ( .A(n12379), .B(n12378), .S(n13053), .Z(n12380) );
  MUX2_X2 U16844 ( .A(decode_regfile_fpregs_18__15_), .B(
        decode_regfile_fpregs_19__15_), .S(n12981), .Z(n12381) );
  MUX2_X2 U16845 ( .A(decode_regfile_fpregs_16__15_), .B(
        decode_regfile_fpregs_17__15_), .S(n12981), .Z(n12382) );
  MUX2_X2 U16846 ( .A(n12382), .B(n12381), .S(n13053), .Z(n12383) );
  MUX2_X2 U16847 ( .A(n12383), .B(n12380), .S(n13078), .Z(n12384) );
  MUX2_X2 U16848 ( .A(n12384), .B(n12377), .S(n13091), .Z(n12385) );
  MUX2_X2 U16849 ( .A(decode_regfile_fpregs_14__15_), .B(
        decode_regfile_fpregs_15__15_), .S(n12982), .Z(n12386) );
  MUX2_X2 U16850 ( .A(decode_regfile_fpregs_12__15_), .B(
        decode_regfile_fpregs_13__15_), .S(n12982), .Z(n12387) );
  MUX2_X2 U16851 ( .A(n12387), .B(n12386), .S(n13054), .Z(n12388) );
  MUX2_X2 U16852 ( .A(decode_regfile_fpregs_10__15_), .B(
        decode_regfile_fpregs_11__15_), .S(n12982), .Z(n12389) );
  MUX2_X2 U16853 ( .A(decode_regfile_fpregs_8__15_), .B(
        decode_regfile_fpregs_9__15_), .S(n12982), .Z(n12390) );
  MUX2_X2 U16854 ( .A(n12390), .B(n12389), .S(n13054), .Z(n12391) );
  MUX2_X2 U16855 ( .A(n12391), .B(n12388), .S(n13079), .Z(n12392) );
  MUX2_X2 U16856 ( .A(decode_regfile_fpregs_6__15_), .B(
        decode_regfile_fpregs_7__15_), .S(n12982), .Z(n12393) );
  MUX2_X2 U16857 ( .A(decode_regfile_fpregs_4__15_), .B(
        decode_regfile_fpregs_5__15_), .S(n12982), .Z(n12394) );
  MUX2_X2 U16858 ( .A(n12394), .B(n12393), .S(n13054), .Z(n12395) );
  MUX2_X2 U16859 ( .A(decode_regfile_fpregs_2__15_), .B(
        decode_regfile_fpregs_3__15_), .S(n12982), .Z(n12396) );
  MUX2_X2 U16860 ( .A(decode_regfile_fpregs_0__15_), .B(
        decode_regfile_fpregs_1__15_), .S(n12982), .Z(n12397) );
  MUX2_X2 U16861 ( .A(n12397), .B(n12396), .S(n13054), .Z(n12398) );
  MUX2_X2 U16862 ( .A(n12398), .B(n12395), .S(n13079), .Z(n12399) );
  MUX2_X2 U16863 ( .A(n12399), .B(n12392), .S(n13092), .Z(n12400) );
  MUX2_X2 U16864 ( .A(n12400), .B(n12385), .S(n13100), .Z(decode_regfile_N148)
         );
  MUX2_X2 U16865 ( .A(decode_regfile_fpregs_30__16_), .B(
        decode_regfile_fpregs_31__16_), .S(n12982), .Z(n12401) );
  MUX2_X2 U16866 ( .A(decode_regfile_fpregs_28__16_), .B(
        decode_regfile_fpregs_29__16_), .S(n12982), .Z(n12402) );
  MUX2_X2 U16867 ( .A(n12402), .B(n12401), .S(n13054), .Z(n12403) );
  MUX2_X2 U16868 ( .A(decode_regfile_fpregs_26__16_), .B(
        decode_regfile_fpregs_27__16_), .S(n12982), .Z(n12404) );
  MUX2_X2 U16869 ( .A(decode_regfile_fpregs_24__16_), .B(
        decode_regfile_fpregs_25__16_), .S(n12983), .Z(n12405) );
  MUX2_X2 U16870 ( .A(n12405), .B(n12404), .S(n13054), .Z(n12406) );
  MUX2_X2 U16871 ( .A(n12406), .B(n12403), .S(n13079), .Z(n12407) );
  MUX2_X2 U16872 ( .A(decode_regfile_fpregs_22__16_), .B(
        decode_regfile_fpregs_23__16_), .S(n12983), .Z(n12408) );
  MUX2_X2 U16873 ( .A(decode_regfile_fpregs_20__16_), .B(
        decode_regfile_fpregs_21__16_), .S(n12983), .Z(n12409) );
  MUX2_X2 U16874 ( .A(n12409), .B(n12408), .S(n13054), .Z(n12410) );
  MUX2_X2 U16875 ( .A(decode_regfile_fpregs_18__16_), .B(
        decode_regfile_fpregs_19__16_), .S(n12983), .Z(n12411) );
  MUX2_X2 U16876 ( .A(decode_regfile_fpregs_16__16_), .B(
        decode_regfile_fpregs_17__16_), .S(n12983), .Z(n12412) );
  MUX2_X2 U16877 ( .A(n12412), .B(n12411), .S(n13054), .Z(n12413) );
  MUX2_X2 U16878 ( .A(n12413), .B(n12410), .S(n13079), .Z(n12414) );
  MUX2_X2 U16879 ( .A(n12414), .B(n12407), .S(n13092), .Z(n12415) );
  MUX2_X2 U16880 ( .A(decode_regfile_fpregs_14__16_), .B(
        decode_regfile_fpregs_15__16_), .S(n12983), .Z(n12416) );
  MUX2_X2 U16881 ( .A(decode_regfile_fpregs_12__16_), .B(
        decode_regfile_fpregs_13__16_), .S(n12983), .Z(n12417) );
  MUX2_X2 U16882 ( .A(n12417), .B(n12416), .S(n13054), .Z(n12418) );
  MUX2_X2 U16883 ( .A(decode_regfile_fpregs_10__16_), .B(
        decode_regfile_fpregs_11__16_), .S(n12983), .Z(n12419) );
  MUX2_X2 U16884 ( .A(decode_regfile_fpregs_8__16_), .B(
        decode_regfile_fpregs_9__16_), .S(n12983), .Z(n12420) );
  MUX2_X2 U16885 ( .A(n12420), .B(n12419), .S(n13054), .Z(n12421) );
  MUX2_X2 U16886 ( .A(n12421), .B(n12418), .S(n13079), .Z(n12422) );
  MUX2_X2 U16887 ( .A(decode_regfile_fpregs_6__16_), .B(
        decode_regfile_fpregs_7__16_), .S(n12983), .Z(n12423) );
  MUX2_X2 U16888 ( .A(decode_regfile_fpregs_4__16_), .B(
        decode_regfile_fpregs_5__16_), .S(n12983), .Z(n12424) );
  MUX2_X2 U16889 ( .A(n12424), .B(n12423), .S(n13054), .Z(n12425) );
  MUX2_X2 U16890 ( .A(decode_regfile_fpregs_2__16_), .B(
        decode_regfile_fpregs_3__16_), .S(n12984), .Z(n12426) );
  MUX2_X2 U16891 ( .A(decode_regfile_fpregs_0__16_), .B(
        decode_regfile_fpregs_1__16_), .S(n12984), .Z(n12427) );
  MUX2_X2 U16892 ( .A(n12427), .B(n12426), .S(n13055), .Z(n12428) );
  MUX2_X2 U16893 ( .A(n12428), .B(n12425), .S(n13079), .Z(n12429) );
  MUX2_X2 U16894 ( .A(n12429), .B(n12422), .S(n13092), .Z(n12430) );
  MUX2_X2 U16895 ( .A(n12430), .B(n12415), .S(n13100), .Z(decode_regfile_N147)
         );
  MUX2_X2 U16896 ( .A(decode_regfile_fpregs_30__17_), .B(
        decode_regfile_fpregs_31__17_), .S(n12984), .Z(n12431) );
  MUX2_X2 U16897 ( .A(decode_regfile_fpregs_28__17_), .B(
        decode_regfile_fpregs_29__17_), .S(n12984), .Z(n12432) );
  MUX2_X2 U16898 ( .A(n12432), .B(n12431), .S(n13055), .Z(n12433) );
  MUX2_X2 U16899 ( .A(decode_regfile_fpregs_26__17_), .B(
        decode_regfile_fpregs_27__17_), .S(n12984), .Z(n12434) );
  MUX2_X2 U16900 ( .A(decode_regfile_fpregs_24__17_), .B(
        decode_regfile_fpregs_25__17_), .S(n12984), .Z(n12435) );
  MUX2_X2 U16901 ( .A(n12435), .B(n12434), .S(n13055), .Z(n12436) );
  MUX2_X2 U16902 ( .A(n12436), .B(n12433), .S(n13079), .Z(n12437) );
  MUX2_X2 U16903 ( .A(decode_regfile_fpregs_22__17_), .B(
        decode_regfile_fpregs_23__17_), .S(n12984), .Z(n12438) );
  MUX2_X2 U16904 ( .A(decode_regfile_fpregs_20__17_), .B(
        decode_regfile_fpregs_21__17_), .S(n12984), .Z(n12439) );
  MUX2_X2 U16905 ( .A(n12439), .B(n12438), .S(n13055), .Z(n12440) );
  MUX2_X2 U16906 ( .A(decode_regfile_fpregs_18__17_), .B(
        decode_regfile_fpregs_19__17_), .S(n12984), .Z(n12441) );
  MUX2_X2 U16907 ( .A(decode_regfile_fpregs_16__17_), .B(
        decode_regfile_fpregs_17__17_), .S(n12984), .Z(n12442) );
  MUX2_X2 U16908 ( .A(n12442), .B(n12441), .S(n13055), .Z(n12443) );
  MUX2_X2 U16909 ( .A(n12443), .B(n12440), .S(n13079), .Z(n12444) );
  MUX2_X2 U16910 ( .A(n12444), .B(n12437), .S(n13092), .Z(n12445) );
  MUX2_X2 U16911 ( .A(decode_regfile_fpregs_14__17_), .B(
        decode_regfile_fpregs_15__17_), .S(n12984), .Z(n12446) );
  MUX2_X2 U16912 ( .A(decode_regfile_fpregs_12__17_), .B(
        decode_regfile_fpregs_13__17_), .S(n12985), .Z(n12447) );
  MUX2_X2 U16913 ( .A(n12447), .B(n12446), .S(n13055), .Z(n12448) );
  MUX2_X2 U16914 ( .A(decode_regfile_fpregs_10__17_), .B(
        decode_regfile_fpregs_11__17_), .S(n12985), .Z(n12449) );
  MUX2_X2 U16915 ( .A(decode_regfile_fpregs_8__17_), .B(
        decode_regfile_fpregs_9__17_), .S(n12985), .Z(n12450) );
  MUX2_X2 U16916 ( .A(n12450), .B(n12449), .S(n13055), .Z(n12451) );
  MUX2_X2 U16917 ( .A(n12451), .B(n12448), .S(n13079), .Z(n12452) );
  MUX2_X2 U16918 ( .A(decode_regfile_fpregs_6__17_), .B(
        decode_regfile_fpregs_7__17_), .S(n12985), .Z(n12453) );
  MUX2_X2 U16919 ( .A(decode_regfile_fpregs_4__17_), .B(
        decode_regfile_fpregs_5__17_), .S(n12985), .Z(n12454) );
  MUX2_X2 U16920 ( .A(n12454), .B(n12453), .S(n13055), .Z(n12455) );
  MUX2_X2 U16921 ( .A(decode_regfile_fpregs_2__17_), .B(
        decode_regfile_fpregs_3__17_), .S(n12985), .Z(n12456) );
  MUX2_X2 U16922 ( .A(decode_regfile_fpregs_0__17_), .B(
        decode_regfile_fpregs_1__17_), .S(n12985), .Z(n12457) );
  MUX2_X2 U16923 ( .A(n12457), .B(n12456), .S(n13055), .Z(n12458) );
  MUX2_X2 U16924 ( .A(n12458), .B(n12455), .S(n13079), .Z(n12459) );
  MUX2_X2 U16925 ( .A(n12459), .B(n12452), .S(n13092), .Z(n12460) );
  MUX2_X2 U16926 ( .A(n12460), .B(n12445), .S(n13100), .Z(decode_regfile_N146)
         );
  MUX2_X2 U16927 ( .A(decode_regfile_fpregs_30__18_), .B(
        decode_regfile_fpregs_31__18_), .S(n12985), .Z(n12461) );
  MUX2_X2 U16928 ( .A(decode_regfile_fpregs_28__18_), .B(
        decode_regfile_fpregs_29__18_), .S(n12985), .Z(n12462) );
  MUX2_X2 U16929 ( .A(n12462), .B(n12461), .S(n13055), .Z(n12463) );
  MUX2_X2 U16930 ( .A(decode_regfile_fpregs_26__18_), .B(
        decode_regfile_fpregs_27__18_), .S(n12985), .Z(n12464) );
  MUX2_X2 U16931 ( .A(decode_regfile_fpregs_24__18_), .B(
        decode_regfile_fpregs_25__18_), .S(n12985), .Z(n12465) );
  MUX2_X2 U16932 ( .A(n12465), .B(n12464), .S(n13055), .Z(n12466) );
  MUX2_X2 U16933 ( .A(n12466), .B(n12463), .S(n13079), .Z(n12467) );
  MUX2_X2 U16934 ( .A(decode_regfile_fpregs_22__18_), .B(
        decode_regfile_fpregs_23__18_), .S(n12986), .Z(n12468) );
  MUX2_X2 U16935 ( .A(decode_regfile_fpregs_20__18_), .B(
        decode_regfile_fpregs_21__18_), .S(n12986), .Z(n12469) );
  MUX2_X2 U16936 ( .A(n12469), .B(n12468), .S(n13056), .Z(n12470) );
  MUX2_X2 U16937 ( .A(decode_regfile_fpregs_18__18_), .B(
        decode_regfile_fpregs_19__18_), .S(n12986), .Z(n12471) );
  MUX2_X2 U16938 ( .A(decode_regfile_fpregs_16__18_), .B(
        decode_regfile_fpregs_17__18_), .S(n12986), .Z(n12472) );
  MUX2_X2 U16939 ( .A(n12472), .B(n12471), .S(n13056), .Z(n12473) );
  MUX2_X2 U16940 ( .A(n12473), .B(n12470), .S(n13080), .Z(n12474) );
  MUX2_X2 U16941 ( .A(n12474), .B(n12467), .S(n13092), .Z(n12475) );
  MUX2_X2 U16942 ( .A(decode_regfile_fpregs_14__18_), .B(
        decode_regfile_fpregs_15__18_), .S(n12986), .Z(n12476) );
  MUX2_X2 U16943 ( .A(decode_regfile_fpregs_12__18_), .B(
        decode_regfile_fpregs_13__18_), .S(n12986), .Z(n12477) );
  MUX2_X2 U16944 ( .A(n12477), .B(n12476), .S(n13056), .Z(n12478) );
  MUX2_X2 U16945 ( .A(decode_regfile_fpregs_10__18_), .B(
        decode_regfile_fpregs_11__18_), .S(n12986), .Z(n12479) );
  MUX2_X2 U16946 ( .A(decode_regfile_fpregs_8__18_), .B(
        decode_regfile_fpregs_9__18_), .S(n12986), .Z(n12480) );
  MUX2_X2 U16947 ( .A(n12480), .B(n12479), .S(n13056), .Z(n12481) );
  MUX2_X2 U16948 ( .A(n12481), .B(n12478), .S(n13080), .Z(n12482) );
  MUX2_X2 U16949 ( .A(decode_regfile_fpregs_6__18_), .B(
        decode_regfile_fpregs_7__18_), .S(n12986), .Z(n12483) );
  MUX2_X2 U16950 ( .A(decode_regfile_fpregs_4__18_), .B(
        decode_regfile_fpregs_5__18_), .S(n12986), .Z(n12484) );
  MUX2_X2 U16951 ( .A(n12484), .B(n12483), .S(n13056), .Z(n12485) );
  MUX2_X2 U16952 ( .A(decode_regfile_fpregs_2__18_), .B(
        decode_regfile_fpregs_3__18_), .S(n12986), .Z(n12486) );
  MUX2_X2 U16953 ( .A(decode_regfile_fpregs_0__18_), .B(
        decode_regfile_fpregs_1__18_), .S(n12987), .Z(n12487) );
  MUX2_X2 U16954 ( .A(n12487), .B(n12486), .S(n13056), .Z(n12488) );
  MUX2_X2 U16955 ( .A(n12488), .B(n12485), .S(n13080), .Z(n12489) );
  MUX2_X2 U16956 ( .A(n12489), .B(n12482), .S(n13092), .Z(n12490) );
  MUX2_X2 U16957 ( .A(n12490), .B(n12475), .S(n13100), .Z(decode_regfile_N145)
         );
  MUX2_X2 U16958 ( .A(decode_regfile_fpregs_30__19_), .B(
        decode_regfile_fpregs_31__19_), .S(n12987), .Z(n12491) );
  MUX2_X2 U16959 ( .A(decode_regfile_fpregs_28__19_), .B(
        decode_regfile_fpregs_29__19_), .S(n12987), .Z(n12492) );
  MUX2_X2 U16960 ( .A(n12492), .B(n12491), .S(n13056), .Z(n12493) );
  MUX2_X2 U16961 ( .A(decode_regfile_fpregs_26__19_), .B(
        decode_regfile_fpregs_27__19_), .S(n12987), .Z(n12494) );
  MUX2_X2 U16962 ( .A(decode_regfile_fpregs_24__19_), .B(
        decode_regfile_fpregs_25__19_), .S(n12987), .Z(n12495) );
  MUX2_X2 U16963 ( .A(n12495), .B(n12494), .S(n13056), .Z(n12496) );
  MUX2_X2 U16964 ( .A(n12496), .B(n12493), .S(n13080), .Z(n12497) );
  MUX2_X2 U16965 ( .A(decode_regfile_fpregs_22__19_), .B(
        decode_regfile_fpregs_23__19_), .S(n12987), .Z(n12498) );
  MUX2_X2 U16966 ( .A(decode_regfile_fpregs_20__19_), .B(
        decode_regfile_fpregs_21__19_), .S(n12987), .Z(n12499) );
  MUX2_X2 U16967 ( .A(n12499), .B(n12498), .S(n13056), .Z(n12500) );
  MUX2_X2 U16968 ( .A(decode_regfile_fpregs_18__19_), .B(
        decode_regfile_fpregs_19__19_), .S(n12987), .Z(n12501) );
  MUX2_X2 U16969 ( .A(decode_regfile_fpregs_16__19_), .B(
        decode_regfile_fpregs_17__19_), .S(n12987), .Z(n12502) );
  MUX2_X2 U16970 ( .A(n12502), .B(n12501), .S(n13056), .Z(n12503) );
  MUX2_X2 U16971 ( .A(n12503), .B(n12500), .S(n13080), .Z(n12504) );
  MUX2_X2 U16972 ( .A(n12504), .B(n12497), .S(n13092), .Z(n12505) );
  MUX2_X2 U16973 ( .A(decode_regfile_fpregs_14__19_), .B(
        decode_regfile_fpregs_15__19_), .S(n12987), .Z(n12506) );
  MUX2_X2 U16974 ( .A(decode_regfile_fpregs_12__19_), .B(
        decode_regfile_fpregs_13__19_), .S(n12987), .Z(n12507) );
  MUX2_X2 U16975 ( .A(n12507), .B(n12506), .S(n13056), .Z(n12508) );
  MUX2_X2 U16976 ( .A(decode_regfile_fpregs_10__19_), .B(
        decode_regfile_fpregs_11__19_), .S(n12988), .Z(n12509) );
  MUX2_X2 U16977 ( .A(decode_regfile_fpregs_8__19_), .B(
        decode_regfile_fpregs_9__19_), .S(n12988), .Z(n12510) );
  MUX2_X2 U16978 ( .A(n12510), .B(n12509), .S(n13015), .Z(n12511) );
  MUX2_X2 U16979 ( .A(n12511), .B(n12508), .S(n13080), .Z(n12512) );
  MUX2_X2 U16980 ( .A(decode_regfile_fpregs_6__19_), .B(
        decode_regfile_fpregs_7__19_), .S(n12988), .Z(n12513) );
  MUX2_X2 U16981 ( .A(decode_regfile_fpregs_4__19_), .B(
        decode_regfile_fpregs_5__19_), .S(n12988), .Z(n12514) );
  MUX2_X2 U16982 ( .A(n12514), .B(n12513), .S(n13009), .Z(n12515) );
  MUX2_X2 U16983 ( .A(decode_regfile_fpregs_2__19_), .B(
        decode_regfile_fpregs_3__19_), .S(n12988), .Z(n12516) );
  MUX2_X2 U16984 ( .A(decode_regfile_fpregs_0__19_), .B(
        decode_regfile_fpregs_1__19_), .S(n12988), .Z(n12517) );
  MUX2_X2 U16985 ( .A(n12517), .B(n12516), .S(n13011), .Z(n12518) );
  MUX2_X2 U16986 ( .A(n12518), .B(n12515), .S(n13080), .Z(n12519) );
  MUX2_X2 U16987 ( .A(n12519), .B(n12512), .S(n13092), .Z(n12520) );
  MUX2_X2 U16988 ( .A(n12520), .B(n12505), .S(n13100), .Z(decode_regfile_N144)
         );
  MUX2_X2 U16989 ( .A(decode_regfile_fpregs_30__20_), .B(
        decode_regfile_fpregs_31__20_), .S(n12988), .Z(n12521) );
  MUX2_X2 U16990 ( .A(decode_regfile_fpregs_28__20_), .B(
        decode_regfile_fpregs_29__20_), .S(n12988), .Z(n12522) );
  MUX2_X2 U16991 ( .A(n12522), .B(n12521), .S(n13008), .Z(n12523) );
  MUX2_X2 U16992 ( .A(decode_regfile_fpregs_26__20_), .B(
        decode_regfile_fpregs_27__20_), .S(n12988), .Z(n12524) );
  MUX2_X2 U16993 ( .A(decode_regfile_fpregs_24__20_), .B(
        decode_regfile_fpregs_25__20_), .S(n12988), .Z(n12525) );
  MUX2_X2 U16994 ( .A(n12525), .B(n12524), .S(n13020), .Z(n12526) );
  MUX2_X2 U16995 ( .A(n12526), .B(n12523), .S(n13080), .Z(n12527) );
  MUX2_X2 U16996 ( .A(decode_regfile_fpregs_22__20_), .B(
        decode_regfile_fpregs_23__20_), .S(n12988), .Z(n12528) );
  MUX2_X2 U16997 ( .A(decode_regfile_fpregs_20__20_), .B(
        decode_regfile_fpregs_21__20_), .S(n12989), .Z(n12529) );
  MUX2_X2 U16998 ( .A(n12529), .B(n12528), .S(n13017), .Z(n12530) );
  MUX2_X2 U16999 ( .A(decode_regfile_fpregs_18__20_), .B(
        decode_regfile_fpregs_19__20_), .S(n12989), .Z(n12531) );
  MUX2_X2 U17000 ( .A(decode_regfile_fpregs_16__20_), .B(
        decode_regfile_fpregs_17__20_), .S(n12989), .Z(n12532) );
  MUX2_X2 U17001 ( .A(n12532), .B(n12531), .S(n13019), .Z(n12533) );
  MUX2_X2 U17002 ( .A(n12533), .B(n12530), .S(n13080), .Z(n12534) );
  MUX2_X2 U17003 ( .A(n12534), .B(n12527), .S(n13092), .Z(n12535) );
  MUX2_X2 U17004 ( .A(decode_regfile_fpregs_14__20_), .B(
        decode_regfile_fpregs_15__20_), .S(n12989), .Z(n12536) );
  MUX2_X2 U17005 ( .A(decode_regfile_fpregs_12__20_), .B(
        decode_regfile_fpregs_13__20_), .S(n12989), .Z(n12537) );
  MUX2_X2 U17006 ( .A(n12537), .B(n12536), .S(n13018), .Z(n12538) );
  MUX2_X2 U17007 ( .A(decode_regfile_fpregs_10__20_), .B(
        decode_regfile_fpregs_11__20_), .S(n12989), .Z(n12539) );
  MUX2_X2 U17008 ( .A(decode_regfile_fpregs_8__20_), .B(
        decode_regfile_fpregs_9__20_), .S(n12989), .Z(n12540) );
  MUX2_X2 U17009 ( .A(n12540), .B(n12539), .S(n13010), .Z(n12541) );
  MUX2_X2 U17010 ( .A(n12541), .B(n12538), .S(n13080), .Z(n12542) );
  MUX2_X2 U17011 ( .A(decode_regfile_fpregs_6__20_), .B(
        decode_regfile_fpregs_7__20_), .S(n12989), .Z(n12543) );
  MUX2_X2 U17012 ( .A(decode_regfile_fpregs_4__20_), .B(
        decode_regfile_fpregs_5__20_), .S(n12989), .Z(n12544) );
  MUX2_X2 U17013 ( .A(n12544), .B(n12543), .S(n13012), .Z(n12545) );
  MUX2_X2 U17014 ( .A(decode_regfile_fpregs_2__20_), .B(
        decode_regfile_fpregs_3__20_), .S(n12989), .Z(n12546) );
  MUX2_X2 U17015 ( .A(decode_regfile_fpregs_0__20_), .B(
        decode_regfile_fpregs_1__20_), .S(n12989), .Z(n12547) );
  MUX2_X2 U17016 ( .A(n12547), .B(n12546), .S(n13008), .Z(n12548) );
  MUX2_X2 U17017 ( .A(n12548), .B(n12545), .S(n13080), .Z(n12549) );
  MUX2_X2 U17018 ( .A(n12549), .B(n12542), .S(n13092), .Z(n12550) );
  MUX2_X2 U17019 ( .A(n12550), .B(n12535), .S(n13100), .Z(decode_regfile_N143)
         );
  MUX2_X2 U17020 ( .A(decode_regfile_fpregs_30__21_), .B(
        decode_regfile_fpregs_31__21_), .S(n12990), .Z(n12551) );
  MUX2_X2 U17021 ( .A(decode_regfile_fpregs_28__21_), .B(
        decode_regfile_fpregs_29__21_), .S(n12990), .Z(n12552) );
  MUX2_X2 U17022 ( .A(n12552), .B(n12551), .S(n13057), .Z(n12553) );
  MUX2_X2 U17023 ( .A(decode_regfile_fpregs_26__21_), .B(
        decode_regfile_fpregs_27__21_), .S(n12990), .Z(n12554) );
  MUX2_X2 U17024 ( .A(decode_regfile_fpregs_24__21_), .B(
        decode_regfile_fpregs_25__21_), .S(n12990), .Z(n12555) );
  MUX2_X2 U17025 ( .A(n12555), .B(n12554), .S(n13057), .Z(n12556) );
  MUX2_X2 U17026 ( .A(n12556), .B(n12553), .S(n13081), .Z(n12557) );
  MUX2_X2 U17027 ( .A(decode_regfile_fpregs_22__21_), .B(
        decode_regfile_fpregs_23__21_), .S(n12990), .Z(n12558) );
  MUX2_X2 U17028 ( .A(decode_regfile_fpregs_20__21_), .B(
        decode_regfile_fpregs_21__21_), .S(n12990), .Z(n12559) );
  MUX2_X2 U17029 ( .A(n12559), .B(n12558), .S(n13057), .Z(n12560) );
  MUX2_X2 U17030 ( .A(decode_regfile_fpregs_18__21_), .B(
        decode_regfile_fpregs_19__21_), .S(n12990), .Z(n12561) );
  MUX2_X2 U17031 ( .A(decode_regfile_fpregs_16__21_), .B(
        decode_regfile_fpregs_17__21_), .S(n12990), .Z(n12562) );
  MUX2_X2 U17032 ( .A(n12562), .B(n12561), .S(n13057), .Z(n12563) );
  MUX2_X2 U17033 ( .A(n12563), .B(n12560), .S(n13081), .Z(n12564) );
  MUX2_X2 U17034 ( .A(n12564), .B(n12557), .S(n13093), .Z(n12565) );
  MUX2_X2 U17035 ( .A(decode_regfile_fpregs_14__21_), .B(
        decode_regfile_fpregs_15__21_), .S(n12990), .Z(n12566) );
  MUX2_X2 U17036 ( .A(decode_regfile_fpregs_12__21_), .B(
        decode_regfile_fpregs_13__21_), .S(n12990), .Z(n12567) );
  MUX2_X2 U17037 ( .A(n12567), .B(n12566), .S(n13057), .Z(n12568) );
  MUX2_X2 U17038 ( .A(decode_regfile_fpregs_10__21_), .B(
        decode_regfile_fpregs_11__21_), .S(n12990), .Z(n12569) );
  MUX2_X2 U17039 ( .A(decode_regfile_fpregs_8__21_), .B(
        decode_regfile_fpregs_9__21_), .S(n12991), .Z(n12570) );
  MUX2_X2 U17040 ( .A(n12570), .B(n12569), .S(n13057), .Z(n12571) );
  MUX2_X2 U17041 ( .A(n12571), .B(n12568), .S(n13081), .Z(n12572) );
  MUX2_X2 U17042 ( .A(decode_regfile_fpregs_6__21_), .B(
        decode_regfile_fpregs_7__21_), .S(n12991), .Z(n12573) );
  MUX2_X2 U17043 ( .A(decode_regfile_fpregs_4__21_), .B(
        decode_regfile_fpregs_5__21_), .S(n12991), .Z(n12574) );
  MUX2_X2 U17044 ( .A(n12574), .B(n12573), .S(n13057), .Z(n12575) );
  MUX2_X2 U17045 ( .A(decode_regfile_fpregs_2__21_), .B(
        decode_regfile_fpregs_3__21_), .S(n12991), .Z(n12576) );
  MUX2_X2 U17046 ( .A(decode_regfile_fpregs_0__21_), .B(
        decode_regfile_fpregs_1__21_), .S(n12991), .Z(n12577) );
  MUX2_X2 U17047 ( .A(n12577), .B(n12576), .S(n13057), .Z(n12578) );
  MUX2_X2 U17048 ( .A(n12578), .B(n12575), .S(n13081), .Z(n12579) );
  MUX2_X2 U17049 ( .A(n12579), .B(n12572), .S(n13093), .Z(n12580) );
  MUX2_X2 U17050 ( .A(n12580), .B(n12565), .S(n13101), .Z(decode_regfile_N142)
         );
  MUX2_X2 U17051 ( .A(decode_regfile_fpregs_30__22_), .B(
        decode_regfile_fpregs_31__22_), .S(n12991), .Z(n12581) );
  MUX2_X2 U17052 ( .A(decode_regfile_fpregs_28__22_), .B(
        decode_regfile_fpregs_29__22_), .S(n12991), .Z(n12582) );
  MUX2_X2 U17053 ( .A(n12582), .B(n12581), .S(n13057), .Z(n12583) );
  MUX2_X2 U17054 ( .A(decode_regfile_fpregs_26__22_), .B(
        decode_regfile_fpregs_27__22_), .S(n12991), .Z(n12584) );
  MUX2_X2 U17055 ( .A(decode_regfile_fpregs_24__22_), .B(
        decode_regfile_fpregs_25__22_), .S(n12991), .Z(n12585) );
  MUX2_X2 U17056 ( .A(n12585), .B(n12584), .S(n13057), .Z(n12586) );
  MUX2_X2 U17057 ( .A(n12586), .B(n12583), .S(n13081), .Z(n12587) );
  MUX2_X2 U17058 ( .A(decode_regfile_fpregs_22__22_), .B(
        decode_regfile_fpregs_23__22_), .S(n12991), .Z(n12588) );
  MUX2_X2 U17059 ( .A(decode_regfile_fpregs_20__22_), .B(
        decode_regfile_fpregs_21__22_), .S(n12991), .Z(n12589) );
  MUX2_X2 U17060 ( .A(n12589), .B(n12588), .S(n13057), .Z(n12590) );
  MUX2_X2 U17061 ( .A(decode_regfile_fpregs_18__22_), .B(
        decode_regfile_fpregs_19__22_), .S(n12992), .Z(n12591) );
  MUX2_X2 U17062 ( .A(decode_regfile_fpregs_16__22_), .B(
        decode_regfile_fpregs_17__22_), .S(n12992), .Z(n12592) );
  MUX2_X2 U17063 ( .A(n12592), .B(n12591), .S(n13058), .Z(n12593) );
  MUX2_X2 U17064 ( .A(n12593), .B(n12590), .S(n13081), .Z(n12594) );
  MUX2_X2 U17065 ( .A(n12594), .B(n12587), .S(n13093), .Z(n12595) );
  MUX2_X2 U17066 ( .A(decode_regfile_fpregs_14__22_), .B(
        decode_regfile_fpregs_15__22_), .S(n12992), .Z(n12596) );
  MUX2_X2 U17067 ( .A(decode_regfile_fpregs_12__22_), .B(
        decode_regfile_fpregs_13__22_), .S(n12992), .Z(n12597) );
  MUX2_X2 U17068 ( .A(n12597), .B(n12596), .S(n13058), .Z(n12598) );
  MUX2_X2 U17069 ( .A(decode_regfile_fpregs_10__22_), .B(
        decode_regfile_fpregs_11__22_), .S(n12992), .Z(n12599) );
  MUX2_X2 U17070 ( .A(decode_regfile_fpregs_8__22_), .B(
        decode_regfile_fpregs_9__22_), .S(n12992), .Z(n12600) );
  MUX2_X2 U17071 ( .A(n12600), .B(n12599), .S(n13058), .Z(n12601) );
  MUX2_X2 U17072 ( .A(n12601), .B(n12598), .S(n13081), .Z(n12602) );
  MUX2_X2 U17073 ( .A(decode_regfile_fpregs_6__22_), .B(
        decode_regfile_fpregs_7__22_), .S(n12992), .Z(n12603) );
  MUX2_X2 U17074 ( .A(decode_regfile_fpregs_4__22_), .B(
        decode_regfile_fpregs_5__22_), .S(n12992), .Z(n12604) );
  MUX2_X2 U17075 ( .A(n12604), .B(n12603), .S(n13058), .Z(n12605) );
  MUX2_X2 U17076 ( .A(decode_regfile_fpregs_2__22_), .B(
        decode_regfile_fpregs_3__22_), .S(n12992), .Z(n12606) );
  MUX2_X2 U17077 ( .A(decode_regfile_fpregs_0__22_), .B(
        decode_regfile_fpregs_1__22_), .S(n12992), .Z(n12607) );
  MUX2_X2 U17078 ( .A(n12607), .B(n12606), .S(n13058), .Z(n12608) );
  MUX2_X2 U17079 ( .A(n12608), .B(n12605), .S(n13081), .Z(n12609) );
  MUX2_X2 U17080 ( .A(n12609), .B(n12602), .S(n13093), .Z(n12610) );
  MUX2_X2 U17081 ( .A(n12610), .B(n12595), .S(n13101), .Z(decode_regfile_N141)
         );
  MUX2_X2 U17082 ( .A(decode_regfile_fpregs_30__23_), .B(
        decode_regfile_fpregs_31__23_), .S(n12992), .Z(n12611) );
  MUX2_X2 U17083 ( .A(decode_regfile_fpregs_28__23_), .B(
        decode_regfile_fpregs_29__23_), .S(n12993), .Z(n12612) );
  MUX2_X2 U17084 ( .A(n12612), .B(n12611), .S(n13058), .Z(n12613) );
  MUX2_X2 U17085 ( .A(decode_regfile_fpregs_26__23_), .B(
        decode_regfile_fpregs_27__23_), .S(n12993), .Z(n12614) );
  MUX2_X2 U17086 ( .A(decode_regfile_fpregs_24__23_), .B(
        decode_regfile_fpregs_25__23_), .S(n12993), .Z(n12615) );
  MUX2_X2 U17087 ( .A(n12615), .B(n12614), .S(n13058), .Z(n12616) );
  MUX2_X2 U17088 ( .A(n12616), .B(n12613), .S(n13081), .Z(n12617) );
  MUX2_X2 U17089 ( .A(decode_regfile_fpregs_22__23_), .B(
        decode_regfile_fpregs_23__23_), .S(n12993), .Z(n12618) );
  MUX2_X2 U17090 ( .A(decode_regfile_fpregs_20__23_), .B(
        decode_regfile_fpregs_21__23_), .S(n12993), .Z(n12619) );
  MUX2_X2 U17091 ( .A(n12619), .B(n12618), .S(n13058), .Z(n12620) );
  MUX2_X2 U17092 ( .A(decode_regfile_fpregs_18__23_), .B(
        decode_regfile_fpregs_19__23_), .S(n12993), .Z(n12621) );
  MUX2_X2 U17093 ( .A(decode_regfile_fpregs_16__23_), .B(
        decode_regfile_fpregs_17__23_), .S(n12993), .Z(n12622) );
  MUX2_X2 U17094 ( .A(n12622), .B(n12621), .S(n13058), .Z(n12623) );
  MUX2_X2 U17095 ( .A(n12623), .B(n12620), .S(n13081), .Z(n12624) );
  MUX2_X2 U17096 ( .A(n12624), .B(n12617), .S(n13093), .Z(n12625) );
  MUX2_X2 U17097 ( .A(decode_regfile_fpregs_14__23_), .B(
        decode_regfile_fpregs_15__23_), .S(n12993), .Z(n12626) );
  MUX2_X2 U17098 ( .A(decode_regfile_fpregs_12__23_), .B(
        decode_regfile_fpregs_13__23_), .S(n12993), .Z(n12627) );
  MUX2_X2 U17099 ( .A(n12627), .B(n12626), .S(n13058), .Z(n12628) );
  MUX2_X2 U17100 ( .A(decode_regfile_fpregs_10__23_), .B(
        decode_regfile_fpregs_11__23_), .S(n12993), .Z(n12629) );
  MUX2_X2 U17101 ( .A(decode_regfile_fpregs_8__23_), .B(
        decode_regfile_fpregs_9__23_), .S(n12993), .Z(n12630) );
  MUX2_X2 U17102 ( .A(n12630), .B(n12629), .S(n13058), .Z(n12631) );
  MUX2_X2 U17103 ( .A(n12631), .B(n12628), .S(n13081), .Z(n12632) );
  MUX2_X2 U17104 ( .A(decode_regfile_fpregs_6__23_), .B(
        decode_regfile_fpregs_7__23_), .S(n12994), .Z(n12633) );
  MUX2_X2 U17105 ( .A(decode_regfile_fpregs_4__23_), .B(
        decode_regfile_fpregs_5__23_), .S(n12994), .Z(n12634) );
  MUX2_X2 U17106 ( .A(n12634), .B(n12633), .S(n13059), .Z(n12635) );
  MUX2_X2 U17107 ( .A(decode_regfile_fpregs_2__23_), .B(
        decode_regfile_fpregs_3__23_), .S(n12994), .Z(n12636) );
  MUX2_X2 U17108 ( .A(decode_regfile_fpregs_0__23_), .B(
        decode_regfile_fpregs_1__23_), .S(n12994), .Z(n12637) );
  MUX2_X2 U17109 ( .A(n12637), .B(n12636), .S(n13059), .Z(n12638) );
  MUX2_X2 U17110 ( .A(n12638), .B(n12635), .S(n13082), .Z(n12639) );
  MUX2_X2 U17111 ( .A(n12639), .B(n12632), .S(n13093), .Z(n12640) );
  MUX2_X2 U17112 ( .A(n12640), .B(n12625), .S(n13101), .Z(decode_regfile_N140)
         );
  MUX2_X2 U17113 ( .A(decode_regfile_fpregs_30__24_), .B(
        decode_regfile_fpregs_31__24_), .S(n12994), .Z(n12641) );
  MUX2_X2 U17114 ( .A(decode_regfile_fpregs_28__24_), .B(
        decode_regfile_fpregs_29__24_), .S(n12994), .Z(n12642) );
  MUX2_X2 U17115 ( .A(n12642), .B(n12641), .S(n13059), .Z(n12643) );
  MUX2_X2 U17116 ( .A(decode_regfile_fpregs_26__24_), .B(
        decode_regfile_fpregs_27__24_), .S(n12994), .Z(n12644) );
  MUX2_X2 U17117 ( .A(decode_regfile_fpregs_24__24_), .B(
        decode_regfile_fpregs_25__24_), .S(n12994), .Z(n12645) );
  MUX2_X2 U17118 ( .A(n12645), .B(n12644), .S(n13059), .Z(n12646) );
  MUX2_X2 U17119 ( .A(n12646), .B(n12643), .S(n13082), .Z(n12647) );
  MUX2_X2 U17120 ( .A(decode_regfile_fpregs_22__24_), .B(
        decode_regfile_fpregs_23__24_), .S(n12994), .Z(n12648) );
  MUX2_X2 U17121 ( .A(decode_regfile_fpregs_20__24_), .B(
        decode_regfile_fpregs_21__24_), .S(n12994), .Z(n12649) );
  MUX2_X2 U17122 ( .A(n12649), .B(n12648), .S(n13059), .Z(n12650) );
  MUX2_X2 U17123 ( .A(decode_regfile_fpregs_18__24_), .B(
        decode_regfile_fpregs_19__24_), .S(n12994), .Z(n12651) );
  MUX2_X2 U17124 ( .A(decode_regfile_fpregs_16__24_), .B(
        decode_regfile_fpregs_17__24_), .S(n12995), .Z(n12652) );
  MUX2_X2 U17125 ( .A(n12652), .B(n12651), .S(n13059), .Z(n12653) );
  MUX2_X2 U17126 ( .A(n12653), .B(n12650), .S(n13082), .Z(n12654) );
  MUX2_X2 U17127 ( .A(n12654), .B(n12647), .S(n13093), .Z(n12655) );
  MUX2_X2 U17128 ( .A(decode_regfile_fpregs_14__24_), .B(
        decode_regfile_fpregs_15__24_), .S(n12995), .Z(n12656) );
  MUX2_X2 U17129 ( .A(decode_regfile_fpregs_12__24_), .B(
        decode_regfile_fpregs_13__24_), .S(n12995), .Z(n12657) );
  MUX2_X2 U17130 ( .A(n12657), .B(n12656), .S(n13059), .Z(n12658) );
  MUX2_X2 U17131 ( .A(decode_regfile_fpregs_10__24_), .B(
        decode_regfile_fpregs_11__24_), .S(n12995), .Z(n12659) );
  MUX2_X2 U17132 ( .A(decode_regfile_fpregs_8__24_), .B(
        decode_regfile_fpregs_9__24_), .S(n12995), .Z(n12660) );
  MUX2_X2 U17133 ( .A(n12660), .B(n12659), .S(n13059), .Z(n12661) );
  MUX2_X2 U17134 ( .A(n12661), .B(n12658), .S(n13082), .Z(n12662) );
  MUX2_X2 U17135 ( .A(decode_regfile_fpregs_6__24_), .B(
        decode_regfile_fpregs_7__24_), .S(n12995), .Z(n12663) );
  MUX2_X2 U17136 ( .A(decode_regfile_fpregs_4__24_), .B(
        decode_regfile_fpregs_5__24_), .S(n12995), .Z(n12664) );
  MUX2_X2 U17137 ( .A(n12664), .B(n12663), .S(n13059), .Z(n12665) );
  MUX2_X2 U17138 ( .A(decode_regfile_fpregs_2__24_), .B(
        decode_regfile_fpregs_3__24_), .S(n12995), .Z(n12666) );
  MUX2_X2 U17139 ( .A(decode_regfile_fpregs_0__24_), .B(
        decode_regfile_fpregs_1__24_), .S(n12995), .Z(n12667) );
  MUX2_X2 U17140 ( .A(n12667), .B(n12666), .S(n13059), .Z(n12668) );
  MUX2_X2 U17141 ( .A(n12668), .B(n12665), .S(n13082), .Z(n12669) );
  MUX2_X2 U17142 ( .A(n12669), .B(n12662), .S(n13093), .Z(n12670) );
  MUX2_X2 U17143 ( .A(n12670), .B(n12655), .S(n13101), .Z(decode_regfile_N139)
         );
  MUX2_X2 U17144 ( .A(decode_regfile_fpregs_30__25_), .B(
        decode_regfile_fpregs_31__25_), .S(n12995), .Z(n12671) );
  MUX2_X2 U17145 ( .A(decode_regfile_fpregs_28__25_), .B(
        decode_regfile_fpregs_29__25_), .S(n12995), .Z(n12672) );
  MUX2_X2 U17146 ( .A(n12672), .B(n12671), .S(n13059), .Z(n12673) );
  MUX2_X2 U17147 ( .A(decode_regfile_fpregs_26__25_), .B(
        decode_regfile_fpregs_27__25_), .S(n12996), .Z(n12674) );
  MUX2_X2 U17148 ( .A(decode_regfile_fpregs_24__25_), .B(
        decode_regfile_fpregs_25__25_), .S(n12996), .Z(n12675) );
  MUX2_X2 U17149 ( .A(n12675), .B(n12674), .S(n13060), .Z(n12676) );
  MUX2_X2 U17150 ( .A(n12676), .B(n12673), .S(n13082), .Z(n12677) );
  MUX2_X2 U17151 ( .A(decode_regfile_fpregs_22__25_), .B(
        decode_regfile_fpregs_23__25_), .S(n12996), .Z(n12678) );
  MUX2_X2 U17152 ( .A(decode_regfile_fpregs_20__25_), .B(
        decode_regfile_fpregs_21__25_), .S(n12996), .Z(n12679) );
  MUX2_X2 U17153 ( .A(n12679), .B(n12678), .S(n13060), .Z(n12680) );
  MUX2_X2 U17154 ( .A(decode_regfile_fpregs_18__25_), .B(
        decode_regfile_fpregs_19__25_), .S(n12996), .Z(n12681) );
  MUX2_X2 U17155 ( .A(decode_regfile_fpregs_16__25_), .B(
        decode_regfile_fpregs_17__25_), .S(n12996), .Z(n12682) );
  MUX2_X2 U17156 ( .A(n12682), .B(n12681), .S(n13060), .Z(n12683) );
  MUX2_X2 U17157 ( .A(n12683), .B(n12680), .S(n13082), .Z(n12684) );
  MUX2_X2 U17158 ( .A(n12684), .B(n12677), .S(n13093), .Z(n12685) );
  MUX2_X2 U17159 ( .A(decode_regfile_fpregs_14__25_), .B(
        decode_regfile_fpregs_15__25_), .S(n12996), .Z(n12686) );
  MUX2_X2 U17160 ( .A(decode_regfile_fpregs_12__25_), .B(
        decode_regfile_fpregs_13__25_), .S(n12996), .Z(n12687) );
  MUX2_X2 U17161 ( .A(n12687), .B(n12686), .S(n13060), .Z(n12688) );
  MUX2_X2 U17162 ( .A(decode_regfile_fpregs_10__25_), .B(
        decode_regfile_fpregs_11__25_), .S(n12996), .Z(n12689) );
  MUX2_X2 U17163 ( .A(decode_regfile_fpregs_8__25_), .B(
        decode_regfile_fpregs_9__25_), .S(n12996), .Z(n12690) );
  MUX2_X2 U17164 ( .A(n12690), .B(n12689), .S(n13060), .Z(n12691) );
  MUX2_X2 U17165 ( .A(n12691), .B(n12688), .S(n13082), .Z(n12692) );
  MUX2_X2 U17166 ( .A(decode_regfile_fpregs_6__25_), .B(
        decode_regfile_fpregs_7__25_), .S(n12996), .Z(n12693) );
  MUX2_X2 U17167 ( .A(decode_regfile_fpregs_4__25_), .B(
        decode_regfile_fpregs_5__25_), .S(n12997), .Z(n12694) );
  MUX2_X2 U17168 ( .A(n12694), .B(n12693), .S(n13060), .Z(n12695) );
  MUX2_X2 U17169 ( .A(decode_regfile_fpregs_2__25_), .B(
        decode_regfile_fpregs_3__25_), .S(n12997), .Z(n12696) );
  MUX2_X2 U17170 ( .A(decode_regfile_fpregs_0__25_), .B(
        decode_regfile_fpregs_1__25_), .S(n12997), .Z(n12697) );
  MUX2_X2 U17171 ( .A(n12697), .B(n12696), .S(n13060), .Z(n12698) );
  MUX2_X2 U17172 ( .A(n12698), .B(n12695), .S(n13082), .Z(n12699) );
  MUX2_X2 U17173 ( .A(n12699), .B(n12692), .S(n13093), .Z(n12700) );
  MUX2_X2 U17174 ( .A(n12700), .B(n12685), .S(n13101), .Z(decode_regfile_N138)
         );
  MUX2_X2 U17175 ( .A(decode_regfile_fpregs_30__26_), .B(
        decode_regfile_fpregs_31__26_), .S(n12997), .Z(n12701) );
  MUX2_X2 U17176 ( .A(decode_regfile_fpregs_28__26_), .B(
        decode_regfile_fpregs_29__26_), .S(n12997), .Z(n12702) );
  MUX2_X2 U17177 ( .A(n12702), .B(n12701), .S(n13060), .Z(n12703) );
  MUX2_X2 U17178 ( .A(decode_regfile_fpregs_26__26_), .B(
        decode_regfile_fpregs_27__26_), .S(n12997), .Z(n12704) );
  MUX2_X2 U17179 ( .A(decode_regfile_fpregs_24__26_), .B(
        decode_regfile_fpregs_25__26_), .S(n12997), .Z(n12705) );
  MUX2_X2 U17180 ( .A(n12705), .B(n12704), .S(n13060), .Z(n12706) );
  MUX2_X2 U17181 ( .A(n12706), .B(n12703), .S(n13082), .Z(n12707) );
  MUX2_X2 U17182 ( .A(decode_regfile_fpregs_22__26_), .B(
        decode_regfile_fpregs_23__26_), .S(n12997), .Z(n12708) );
  MUX2_X2 U17183 ( .A(decode_regfile_fpregs_20__26_), .B(
        decode_regfile_fpregs_21__26_), .S(n12997), .Z(n12709) );
  MUX2_X2 U17184 ( .A(n12709), .B(n12708), .S(n13060), .Z(n12710) );
  MUX2_X2 U17185 ( .A(decode_regfile_fpregs_18__26_), .B(
        decode_regfile_fpregs_19__26_), .S(n12997), .Z(n12711) );
  MUX2_X2 U17186 ( .A(decode_regfile_fpregs_16__26_), .B(
        decode_regfile_fpregs_17__26_), .S(n12997), .Z(n12712) );
  MUX2_X2 U17187 ( .A(n12712), .B(n12711), .S(n13060), .Z(n12713) );
  MUX2_X2 U17188 ( .A(n12713), .B(n12710), .S(n13082), .Z(n12714) );
  MUX2_X2 U17189 ( .A(n12714), .B(n12707), .S(n13093), .Z(n12715) );
  MUX2_X2 U17190 ( .A(decode_regfile_fpregs_14__26_), .B(
        decode_regfile_fpregs_15__26_), .S(n12998), .Z(n12716) );
  MUX2_X2 U17191 ( .A(decode_regfile_fpregs_12__26_), .B(
        decode_regfile_fpregs_13__26_), .S(n12998), .Z(n12717) );
  MUX2_X2 U17192 ( .A(n12717), .B(n12716), .S(n13018), .Z(n12718) );
  MUX2_X2 U17193 ( .A(decode_regfile_fpregs_10__26_), .B(
        decode_regfile_fpregs_11__26_), .S(n12998), .Z(n12719) );
  MUX2_X2 U17194 ( .A(decode_regfile_fpregs_8__26_), .B(
        decode_regfile_fpregs_9__26_), .S(n12998), .Z(n12720) );
  MUX2_X2 U17195 ( .A(n12720), .B(n12719), .S(n13012), .Z(n12721) );
  MUX2_X2 U17196 ( .A(n12721), .B(n12718), .S(n13083), .Z(n12722) );
  MUX2_X2 U17197 ( .A(decode_regfile_fpregs_6__26_), .B(
        decode_regfile_fpregs_7__26_), .S(n12998), .Z(n12723) );
  MUX2_X2 U17198 ( .A(decode_regfile_fpregs_4__26_), .B(
        decode_regfile_fpregs_5__26_), .S(n12998), .Z(n12724) );
  MUX2_X2 U17199 ( .A(n12724), .B(n12723), .S(n13011), .Z(n12725) );
  MUX2_X2 U17200 ( .A(decode_regfile_fpregs_2__26_), .B(
        decode_regfile_fpregs_3__26_), .S(n12998), .Z(n12726) );
  MUX2_X2 U17201 ( .A(decode_regfile_fpregs_0__26_), .B(
        decode_regfile_fpregs_1__26_), .S(n12998), .Z(n12727) );
  MUX2_X2 U17202 ( .A(n12727), .B(n12726), .S(n13006), .Z(n12728) );
  MUX2_X2 U17203 ( .A(n12728), .B(n12725), .S(n13083), .Z(n12729) );
  MUX2_X2 U17204 ( .A(n12729), .B(n12722), .S(n13094), .Z(n12730) );
  MUX2_X2 U17205 ( .A(n12730), .B(n12715), .S(n13101), .Z(decode_regfile_N137)
         );
  MUX2_X2 U17206 ( .A(decode_regfile_fpregs_30__27_), .B(
        decode_regfile_fpregs_31__27_), .S(n12998), .Z(n12731) );
  MUX2_X2 U17207 ( .A(decode_regfile_fpregs_28__27_), .B(
        decode_regfile_fpregs_29__27_), .S(n12998), .Z(n12732) );
  MUX2_X2 U17208 ( .A(n12732), .B(n12731), .S(n13006), .Z(n12733) );
  MUX2_X2 U17209 ( .A(decode_regfile_fpregs_26__27_), .B(
        decode_regfile_fpregs_27__27_), .S(n12998), .Z(n12734) );
  MUX2_X2 U17210 ( .A(decode_regfile_fpregs_24__27_), .B(
        decode_regfile_fpregs_25__27_), .S(n12999), .Z(n12735) );
  MUX2_X2 U17211 ( .A(n12735), .B(n12734), .S(n13019), .Z(n12736) );
  MUX2_X2 U17212 ( .A(n12736), .B(n12733), .S(n13083), .Z(n12737) );
  MUX2_X2 U17213 ( .A(decode_regfile_fpregs_22__27_), .B(
        decode_regfile_fpregs_23__27_), .S(n12999), .Z(n12738) );
  MUX2_X2 U17214 ( .A(decode_regfile_fpregs_20__27_), .B(
        decode_regfile_fpregs_21__27_), .S(n12999), .Z(n12739) );
  MUX2_X2 U17215 ( .A(n12739), .B(n12738), .S(n13017), .Z(n12740) );
  MUX2_X2 U17216 ( .A(decode_regfile_fpregs_18__27_), .B(
        decode_regfile_fpregs_19__27_), .S(n12999), .Z(n12741) );
  MUX2_X2 U17217 ( .A(decode_regfile_fpregs_16__27_), .B(
        decode_regfile_fpregs_17__27_), .S(n12999), .Z(n12742) );
  MUX2_X2 U17218 ( .A(n12742), .B(n12741), .S(n13009), .Z(n12743) );
  MUX2_X2 U17219 ( .A(n12743), .B(n12740), .S(n13083), .Z(n12744) );
  MUX2_X2 U17220 ( .A(n12744), .B(n12737), .S(n13094), .Z(n12745) );
  MUX2_X2 U17221 ( .A(decode_regfile_fpregs_14__27_), .B(
        decode_regfile_fpregs_15__27_), .S(n12999), .Z(n12746) );
  MUX2_X2 U17222 ( .A(decode_regfile_fpregs_12__27_), .B(
        decode_regfile_fpregs_13__27_), .S(n12999), .Z(n12747) );
  MUX2_X2 U17223 ( .A(n12747), .B(n12746), .S(n13015), .Z(n12748) );
  MUX2_X2 U17224 ( .A(decode_regfile_fpregs_10__27_), .B(
        decode_regfile_fpregs_11__27_), .S(n12999), .Z(n12749) );
  MUX2_X2 U17225 ( .A(decode_regfile_fpregs_8__27_), .B(
        decode_regfile_fpregs_9__27_), .S(n12999), .Z(n12750) );
  MUX2_X2 U17226 ( .A(n12750), .B(n12749), .S(n13008), .Z(n12751) );
  MUX2_X2 U17227 ( .A(n12751), .B(n12748), .S(n13083), .Z(n12752) );
  MUX2_X2 U17228 ( .A(decode_regfile_fpregs_6__27_), .B(
        decode_regfile_fpregs_7__27_), .S(n12999), .Z(n12753) );
  MUX2_X2 U17229 ( .A(decode_regfile_fpregs_4__27_), .B(
        decode_regfile_fpregs_5__27_), .S(n12999), .Z(n12754) );
  MUX2_X2 U17230 ( .A(n12754), .B(n12753), .S(n13010), .Z(n12755) );
  MUX2_X2 U17231 ( .A(decode_regfile_fpregs_2__27_), .B(
        decode_regfile_fpregs_3__27_), .S(n13000), .Z(n12756) );
  MUX2_X2 U17232 ( .A(decode_regfile_fpregs_0__27_), .B(
        decode_regfile_fpregs_1__27_), .S(n13000), .Z(n12757) );
  MUX2_X2 U17233 ( .A(n12757), .B(n12756), .S(n13015), .Z(n12758) );
  MUX2_X2 U17234 ( .A(n12758), .B(n12755), .S(n13083), .Z(n12759) );
  MUX2_X2 U17235 ( .A(n12759), .B(n12752), .S(n13094), .Z(n12760) );
  MUX2_X2 U17236 ( .A(n12760), .B(n12745), .S(n13101), .Z(decode_regfile_N136)
         );
  MUX2_X2 U17237 ( .A(decode_regfile_fpregs_30__28_), .B(
        decode_regfile_fpregs_31__28_), .S(n13000), .Z(n12761) );
  MUX2_X2 U17238 ( .A(decode_regfile_fpregs_28__28_), .B(
        decode_regfile_fpregs_29__28_), .S(n13000), .Z(n12762) );
  MUX2_X2 U17239 ( .A(n12762), .B(n12761), .S(n13006), .Z(n12763) );
  MUX2_X2 U17240 ( .A(decode_regfile_fpregs_26__28_), .B(
        decode_regfile_fpregs_27__28_), .S(n13000), .Z(n12764) );
  MUX2_X2 U17241 ( .A(decode_regfile_fpregs_24__28_), .B(
        decode_regfile_fpregs_25__28_), .S(n13000), .Z(n12765) );
  MUX2_X2 U17242 ( .A(n12765), .B(n12764), .S(n13007), .Z(n12766) );
  MUX2_X2 U17243 ( .A(n12766), .B(n12763), .S(n13083), .Z(n12767) );
  MUX2_X2 U17244 ( .A(decode_regfile_fpregs_22__28_), .B(
        decode_regfile_fpregs_23__28_), .S(n13000), .Z(n12768) );
  MUX2_X2 U17245 ( .A(decode_regfile_fpregs_20__28_), .B(
        decode_regfile_fpregs_21__28_), .S(n13000), .Z(n12769) );
  MUX2_X2 U17246 ( .A(n12769), .B(n12768), .S(n13013), .Z(n12770) );
  MUX2_X2 U17247 ( .A(decode_regfile_fpregs_18__28_), .B(
        decode_regfile_fpregs_19__28_), .S(n13000), .Z(n12771) );
  MUX2_X2 U17248 ( .A(decode_regfile_fpregs_16__28_), .B(
        decode_regfile_fpregs_17__28_), .S(n13000), .Z(n12772) );
  MUX2_X2 U17249 ( .A(n12772), .B(n12771), .S(n13017), .Z(n12773) );
  MUX2_X2 U17250 ( .A(n12773), .B(n12770), .S(n13083), .Z(n12774) );
  MUX2_X2 U17251 ( .A(n12774), .B(n12767), .S(n13094), .Z(n12775) );
  MUX2_X2 U17252 ( .A(decode_regfile_fpregs_14__28_), .B(
        decode_regfile_fpregs_15__28_), .S(n13000), .Z(n12776) );
  MUX2_X2 U17253 ( .A(decode_regfile_fpregs_12__28_), .B(
        decode_regfile_fpregs_13__28_), .S(n13001), .Z(n12777) );
  MUX2_X2 U17254 ( .A(n12777), .B(n12776), .S(n13016), .Z(n12778) );
  MUX2_X2 U17255 ( .A(decode_regfile_fpregs_10__28_), .B(
        decode_regfile_fpregs_11__28_), .S(n13001), .Z(n12779) );
  MUX2_X2 U17256 ( .A(decode_regfile_fpregs_8__28_), .B(
        decode_regfile_fpregs_9__28_), .S(n13001), .Z(n12780) );
  MUX2_X2 U17257 ( .A(n12780), .B(n12779), .S(n13018), .Z(n12781) );
  MUX2_X2 U17258 ( .A(n12781), .B(n12778), .S(n13083), .Z(n12782) );
  MUX2_X2 U17259 ( .A(decode_regfile_fpregs_6__28_), .B(
        decode_regfile_fpregs_7__28_), .S(n13001), .Z(n12783) );
  MUX2_X2 U17260 ( .A(decode_regfile_fpregs_4__28_), .B(
        decode_regfile_fpregs_5__28_), .S(n13001), .Z(n12784) );
  MUX2_X2 U17261 ( .A(n12784), .B(n12783), .S(n13019), .Z(n12785) );
  MUX2_X2 U17262 ( .A(decode_regfile_fpregs_2__28_), .B(
        decode_regfile_fpregs_3__28_), .S(n13001), .Z(n12786) );
  MUX2_X2 U17263 ( .A(decode_regfile_fpregs_0__28_), .B(
        decode_regfile_fpregs_1__28_), .S(n13001), .Z(n12787) );
  MUX2_X2 U17264 ( .A(n12787), .B(n12786), .S(n13009), .Z(n12788) );
  MUX2_X2 U17265 ( .A(n12788), .B(n12785), .S(n13083), .Z(n12789) );
  MUX2_X2 U17266 ( .A(n12789), .B(n12782), .S(n13094), .Z(n12790) );
  MUX2_X2 U17267 ( .A(n12790), .B(n12775), .S(n13101), .Z(decode_regfile_N135)
         );
  MUX2_X2 U17268 ( .A(decode_regfile_fpregs_30__29_), .B(
        decode_regfile_fpregs_31__29_), .S(n13001), .Z(n12791) );
  MUX2_X2 U17269 ( .A(decode_regfile_fpregs_28__29_), .B(
        decode_regfile_fpregs_29__29_), .S(n13001), .Z(n12792) );
  MUX2_X2 U17270 ( .A(n12792), .B(n12791), .S(n13014), .Z(n12793) );
  MUX2_X2 U17271 ( .A(decode_regfile_fpregs_26__29_), .B(
        decode_regfile_fpregs_27__29_), .S(n13001), .Z(n12794) );
  MUX2_X2 U17272 ( .A(decode_regfile_fpregs_24__29_), .B(
        decode_regfile_fpregs_25__29_), .S(n13001), .Z(n12795) );
  MUX2_X2 U17273 ( .A(n12795), .B(n12794), .S(n13020), .Z(n12796) );
  MUX2_X2 U17274 ( .A(n12796), .B(n12793), .S(n13083), .Z(n12797) );
  MUX2_X2 U17275 ( .A(decode_regfile_fpregs_22__29_), .B(
        decode_regfile_fpregs_23__29_), .S(n13002), .Z(n12798) );
  MUX2_X2 U17276 ( .A(decode_regfile_fpregs_20__29_), .B(
        decode_regfile_fpregs_21__29_), .S(n13002), .Z(n12799) );
  MUX2_X2 U17277 ( .A(n12799), .B(n12798), .S(n13005), .Z(n12800) );
  MUX2_X2 U17278 ( .A(decode_regfile_fpregs_18__29_), .B(
        decode_regfile_fpregs_19__29_), .S(n13002), .Z(n12801) );
  MUX2_X2 U17279 ( .A(decode_regfile_fpregs_16__29_), .B(
        decode_regfile_fpregs_17__29_), .S(n13002), .Z(n12802) );
  MUX2_X2 U17280 ( .A(n12802), .B(n12801), .S(n13005), .Z(n12803) );
  MUX2_X2 U17281 ( .A(n12803), .B(n12800), .S(n13061), .Z(n12804) );
  MUX2_X2 U17282 ( .A(n12804), .B(n12797), .S(n13094), .Z(n12805) );
  MUX2_X2 U17283 ( .A(decode_regfile_fpregs_14__29_), .B(
        decode_regfile_fpregs_15__29_), .S(n13002), .Z(n12806) );
  MUX2_X2 U17284 ( .A(decode_regfile_fpregs_12__29_), .B(
        decode_regfile_fpregs_13__29_), .S(n13002), .Z(n12807) );
  MUX2_X2 U17285 ( .A(n12807), .B(n12806), .S(n13005), .Z(n12808) );
  MUX2_X2 U17286 ( .A(decode_regfile_fpregs_10__29_), .B(
        decode_regfile_fpregs_11__29_), .S(n13002), .Z(n12809) );
  MUX2_X2 U17287 ( .A(decode_regfile_fpregs_8__29_), .B(
        decode_regfile_fpregs_9__29_), .S(n13002), .Z(n12810) );
  MUX2_X2 U17288 ( .A(n12810), .B(n12809), .S(n13005), .Z(n12811) );
  MUX2_X2 U17289 ( .A(n12811), .B(n12808), .S(n13061), .Z(n12812) );
  MUX2_X2 U17290 ( .A(decode_regfile_fpregs_6__29_), .B(
        decode_regfile_fpregs_7__29_), .S(n13002), .Z(n12813) );
  MUX2_X2 U17291 ( .A(decode_regfile_fpregs_4__29_), .B(
        decode_regfile_fpregs_5__29_), .S(n13002), .Z(n12814) );
  MUX2_X2 U17292 ( .A(n12814), .B(n12813), .S(n13005), .Z(n12815) );
  MUX2_X2 U17293 ( .A(decode_regfile_fpregs_2__29_), .B(
        decode_regfile_fpregs_3__29_), .S(n13002), .Z(n12816) );
  MUX2_X2 U17294 ( .A(decode_regfile_fpregs_0__29_), .B(
        decode_regfile_fpregs_1__29_), .S(n13003), .Z(n12817) );
  MUX2_X2 U17295 ( .A(n12817), .B(n12816), .S(n13011), .Z(n12818) );
  MUX2_X2 U17296 ( .A(n12818), .B(n12815), .S(n13078), .Z(n12819) );
  MUX2_X2 U17297 ( .A(n12819), .B(n12812), .S(n13094), .Z(n12820) );
  MUX2_X2 U17298 ( .A(n12820), .B(n12805), .S(n13101), .Z(decode_regfile_N134)
         );
  MUX2_X2 U17299 ( .A(decode_regfile_fpregs_30__30_), .B(
        decode_regfile_fpregs_31__30_), .S(n13003), .Z(n12821) );
  MUX2_X2 U17300 ( .A(decode_regfile_fpregs_28__30_), .B(
        decode_regfile_fpregs_29__30_), .S(n13003), .Z(n12822) );
  MUX2_X2 U17301 ( .A(n12822), .B(n12821), .S(n13005), .Z(n12823) );
  MUX2_X2 U17302 ( .A(decode_regfile_fpregs_26__30_), .B(
        decode_regfile_fpregs_27__30_), .S(n13003), .Z(n12824) );
  MUX2_X2 U17303 ( .A(decode_regfile_fpregs_24__30_), .B(
        decode_regfile_fpregs_25__30_), .S(n13003), .Z(n12825) );
  MUX2_X2 U17304 ( .A(n12825), .B(n12824), .S(n13005), .Z(n12826) );
  MUX2_X2 U17305 ( .A(n12826), .B(n12823), .S(n13061), .Z(n12827) );
  MUX2_X2 U17306 ( .A(decode_regfile_fpregs_22__30_), .B(
        decode_regfile_fpregs_23__30_), .S(n13003), .Z(n12828) );
  MUX2_X2 U17307 ( .A(decode_regfile_fpregs_20__30_), .B(
        decode_regfile_fpregs_21__30_), .S(n13003), .Z(n12829) );
  MUX2_X2 U17308 ( .A(n12829), .B(n12828), .S(n13005), .Z(n12830) );
  MUX2_X2 U17309 ( .A(decode_regfile_fpregs_18__30_), .B(
        decode_regfile_fpregs_19__30_), .S(n13003), .Z(n12831) );
  MUX2_X2 U17310 ( .A(decode_regfile_fpregs_16__30_), .B(
        decode_regfile_fpregs_17__30_), .S(n13003), .Z(n12832) );
  MUX2_X2 U17311 ( .A(n12832), .B(n12831), .S(n13005), .Z(n12833) );
  MUX2_X2 U17312 ( .A(n12833), .B(n12830), .S(n13061), .Z(n12834) );
  MUX2_X2 U17313 ( .A(n12834), .B(n12827), .S(n13094), .Z(n12835) );
  MUX2_X2 U17314 ( .A(decode_regfile_fpregs_14__30_), .B(
        decode_regfile_fpregs_15__30_), .S(n13003), .Z(n12836) );
  MUX2_X2 U17315 ( .A(decode_regfile_fpregs_12__30_), .B(
        decode_regfile_fpregs_13__30_), .S(n13003), .Z(n12837) );
  MUX2_X2 U17316 ( .A(n12837), .B(n12836), .S(n13005), .Z(n12838) );
  MUX2_X2 U17317 ( .A(decode_regfile_fpregs_10__30_), .B(
        decode_regfile_fpregs_11__30_), .S(n13004), .Z(n12839) );
  MUX2_X2 U17318 ( .A(decode_regfile_fpregs_8__30_), .B(
        decode_regfile_fpregs_9__30_), .S(n13004), .Z(n12840) );
  MUX2_X2 U17319 ( .A(n12840), .B(n12839), .S(n13021), .Z(n12841) );
  MUX2_X2 U17320 ( .A(n12841), .B(n12838), .S(n13061), .Z(n12842) );
  MUX2_X2 U17321 ( .A(decode_regfile_fpregs_6__30_), .B(
        decode_regfile_fpregs_7__30_), .S(n13004), .Z(n12843) );
  MUX2_X2 U17322 ( .A(decode_regfile_fpregs_4__30_), .B(
        decode_regfile_fpregs_5__30_), .S(n13004), .Z(n12844) );
  MUX2_X2 U17323 ( .A(n12844), .B(n12843), .S(n13014), .Z(n12845) );
  MUX2_X2 U17324 ( .A(decode_regfile_fpregs_2__30_), .B(
        decode_regfile_fpregs_3__30_), .S(n13004), .Z(n12846) );
  MUX2_X2 U17325 ( .A(decode_regfile_fpregs_0__30_), .B(
        decode_regfile_fpregs_1__30_), .S(n13004), .Z(n12847) );
  MUX2_X2 U17326 ( .A(n12847), .B(n12846), .S(n13013), .Z(n12848) );
  MUX2_X2 U17327 ( .A(n12848), .B(n12845), .S(n13077), .Z(n12849) );
  MUX2_X2 U17328 ( .A(n12849), .B(n12842), .S(n13094), .Z(n12850) );
  MUX2_X2 U17329 ( .A(n12850), .B(n12835), .S(n13101), .Z(decode_regfile_N133)
         );
  MUX2_X2 U17330 ( .A(decode_regfile_fpregs_30__31_), .B(
        decode_regfile_fpregs_31__31_), .S(n13004), .Z(n12851) );
  MUX2_X2 U17331 ( .A(decode_regfile_fpregs_28__31_), .B(
        decode_regfile_fpregs_29__31_), .S(n13004), .Z(n12852) );
  MUX2_X2 U17332 ( .A(n12852), .B(n12851), .S(n13005), .Z(n12853) );
  MUX2_X2 U17333 ( .A(decode_regfile_fpregs_26__31_), .B(
        decode_regfile_fpregs_27__31_), .S(n13004), .Z(n12854) );
  MUX2_X2 U17334 ( .A(decode_regfile_fpregs_24__31_), .B(
        decode_regfile_fpregs_25__31_), .S(n13004), .Z(n12855) );
  MUX2_X2 U17335 ( .A(n12855), .B(n12854), .S(n13005), .Z(n12856) );
  MUX2_X2 U17336 ( .A(n12856), .B(n12853), .S(n13061), .Z(n12857) );
  MUX2_X2 U17337 ( .A(decode_regfile_fpregs_22__31_), .B(
        decode_regfile_fpregs_23__31_), .S(n13004), .Z(n12858) );
  MUX2_X2 U17338 ( .A(decode_regfile_fpregs_20__31_), .B(
        decode_regfile_fpregs_21__31_), .S(n12881), .Z(n12859) );
  MUX2_X2 U17339 ( .A(n12859), .B(n12858), .S(n13021), .Z(n12860) );
  MUX2_X2 U17340 ( .A(decode_regfile_fpregs_18__31_), .B(
        decode_regfile_fpregs_19__31_), .S(n12912), .Z(n12861) );
  MUX2_X2 U17341 ( .A(decode_regfile_fpregs_16__31_), .B(
        decode_regfile_fpregs_17__31_), .S(n12881), .Z(n12862) );
  MUX2_X2 U17342 ( .A(n12862), .B(n12861), .S(n13021), .Z(n12863) );
  MUX2_X2 U17343 ( .A(n12863), .B(n12860), .S(n13061), .Z(n12864) );
  MUX2_X2 U17344 ( .A(n12864), .B(n12857), .S(n13094), .Z(n12865) );
  MUX2_X2 U17345 ( .A(decode_regfile_fpregs_14__31_), .B(
        decode_regfile_fpregs_15__31_), .S(n12881), .Z(n12866) );
  MUX2_X2 U17346 ( .A(decode_regfile_fpregs_12__31_), .B(
        decode_regfile_fpregs_13__31_), .S(n12881), .Z(n12867) );
  MUX2_X2 U17347 ( .A(n12867), .B(n12866), .S(n13021), .Z(n12868) );
  MUX2_X2 U17348 ( .A(decode_regfile_fpregs_10__31_), .B(
        decode_regfile_fpregs_11__31_), .S(n12881), .Z(n12869) );
  MUX2_X2 U17349 ( .A(decode_regfile_fpregs_8__31_), .B(
        decode_regfile_fpregs_9__31_), .S(n12881), .Z(n12870) );
  MUX2_X2 U17350 ( .A(n12870), .B(n12869), .S(n13007), .Z(n12871) );
  MUX2_X2 U17351 ( .A(n12871), .B(n12868), .S(n13061), .Z(n12872) );
  MUX2_X2 U17352 ( .A(decode_regfile_fpregs_6__31_), .B(
        decode_regfile_fpregs_7__31_), .S(n12881), .Z(n12873) );
  MUX2_X2 U17353 ( .A(decode_regfile_fpregs_4__31_), .B(
        decode_regfile_fpregs_5__31_), .S(n12881), .Z(n12874) );
  MUX2_X2 U17354 ( .A(n12874), .B(n12873), .S(n13006), .Z(n12875) );
  MUX2_X2 U17355 ( .A(decode_regfile_fpregs_2__31_), .B(
        decode_regfile_fpregs_3__31_), .S(n12881), .Z(n12876) );
  MUX2_X2 U17356 ( .A(decode_regfile_fpregs_0__31_), .B(
        decode_regfile_fpregs_1__31_), .S(n12881), .Z(n12877) );
  MUX2_X2 U17357 ( .A(n12877), .B(n12876), .S(n13016), .Z(n12878) );
  MUX2_X2 U17358 ( .A(n12878), .B(n12875), .S(n13076), .Z(n12879) );
  MUX2_X2 U17359 ( .A(n12879), .B(n12872), .S(n13094), .Z(n12880) );
  MUX2_X2 U17360 ( .A(n12880), .B(n12865), .S(n13101), .Z(decode_regfile_N132)
         );
  AND2_X4 U17361 ( .A1(n5358), .A2(n16469), .ZN(n2726) );
  AND2_X4 U17362 ( .A1(n5358), .A2(n8696), .ZN(n2724) );
  AND2_X4 U17363 ( .A1(rw_3[1]), .A2(n8754), .ZN(n733) );
  AND2_X4 U17364 ( .A1(rw_3[1]), .A2(rw_3[0]), .ZN(n699) );
  NOR2_X1 U17365 ( .A1(n13802), .A2(rw_3[0]), .ZN(n13810) );
  OAI22_X1 U17366 ( .A1(n13810), .A2(n8755), .B1(decode_rs2_1_), .B2(n13810), 
        .ZN(n13814) );
  AND2_X1 U17367 ( .A1(rw_3[0]), .A2(n13802), .ZN(n13811) );
  OAI22_X1 U17368 ( .A1(rw_3[1]), .A2(n13811), .B1(n13811), .B2(n13800), .ZN(
        n13813) );
  XNOR2_X1 U17369 ( .A(n13798), .B(rw_3[2]), .ZN(n13812) );
  NAND3_X1 U17370 ( .A1(n13814), .A2(n13813), .A3(n13812), .ZN(n13817) );
  XOR2_X1 U17371 ( .A(decode_rs2_3_), .B(rw_3[3]), .Z(n13816) );
  XOR2_X1 U17372 ( .A(decode_rs2_4_), .B(rw_3[4]), .Z(n13815) );
  NOR3_X1 U17373 ( .A1(n13817), .A2(n13816), .A3(n13815), .ZN(decode_N4) );
  NOR2_X1 U17374 ( .A1(n8810), .A2(rw_3[0]), .ZN(n13818) );
  OAI22_X1 U17375 ( .A1(n13818), .A2(n8755), .B1(n13796), .B2(n13818), .ZN(
        n13822) );
  AND2_X1 U17376 ( .A1(rw_3[0]), .A2(n8810), .ZN(n13819) );
  OAI22_X1 U17377 ( .A1(rw_3[1]), .A2(n13819), .B1(n13819), .B2(n8811), .ZN(
        n13821) );
  XNOR2_X1 U17378 ( .A(decode_rs1_2_), .B(rw_3[2]), .ZN(n13820) );
  NAND3_X1 U17379 ( .A1(n13822), .A2(n13821), .A3(n13820), .ZN(n13825) );
  XOR2_X1 U17380 ( .A(decode_rs1_3_), .B(rw_3[3]), .Z(n13824) );
  XOR2_X1 U17381 ( .A(decode_rs1_4_), .B(rw_3[4]), .Z(n13823) );
  NOR3_X1 U17382 ( .A1(n13825), .A2(n13824), .A3(n13823), .ZN(decode_N2) );
  NOR2_X1 U17383 ( .A1(n8803), .A2(instruction_1[16]), .ZN(n13826) );
  OAI22_X1 U17384 ( .A1(n13826), .A2(n8804), .B1(rw_2[1]), .B2(n13826), .ZN(
        n13830) );
  AND2_X1 U17385 ( .A1(instruction_1[16]), .A2(n8803), .ZN(n13827) );
  OAI22_X1 U17386 ( .A1(instruction_1[17]), .A2(n13827), .B1(n13827), .B2(
        n8806), .ZN(n13829) );
  XNOR2_X1 U17387 ( .A(rw_2[2]), .B(instruction_1[18]), .ZN(n13828) );
  NAND3_X1 U17388 ( .A1(n13830), .A2(n13829), .A3(n13828), .ZN(n13833) );
  XOR2_X1 U17389 ( .A(rw_2[3]), .B(instruction_1[19]), .Z(n13832) );
  XOR2_X1 U17390 ( .A(rw_2[4]), .B(instruction_1[20]), .Z(n13831) );
  NOR3_X1 U17391 ( .A1(n13833), .A2(n13832), .A3(n13831), .ZN(N34) );
  NOR2_X1 U17392 ( .A1(n8795), .A2(instruction_1[16]), .ZN(n13834) );
  OAI22_X1 U17393 ( .A1(n13834), .A2(n8804), .B1(rw_1[1]), .B2(n13834), .ZN(
        n13838) );
  AND2_X1 U17394 ( .A1(instruction_1[16]), .A2(n8795), .ZN(n13835) );
  OAI22_X1 U17395 ( .A1(instruction_1[17]), .A2(n13835), .B1(n13835), .B2(
        n8796), .ZN(n13837) );
  XNOR2_X1 U17396 ( .A(rw_1[2]), .B(instruction_1[18]), .ZN(n13836) );
  NAND3_X1 U17397 ( .A1(n13838), .A2(n13837), .A3(n13836), .ZN(n13841) );
  XOR2_X1 U17398 ( .A(rw_1[3]), .B(instruction_1[19]), .Z(n13840) );
  XOR2_X1 U17399 ( .A(rw_1[4]), .B(instruction_1[20]), .Z(n13839) );
  NOR3_X1 U17400 ( .A1(n13841), .A2(n13840), .A3(n13839), .ZN(N32) );
  NOR2_X1 U17401 ( .A1(n8803), .A2(instruction_1[21]), .ZN(n13842) );
  OAI22_X1 U17402 ( .A1(n13842), .A2(n8805), .B1(rw_2[1]), .B2(n13842), .ZN(
        n13846) );
  AND2_X1 U17403 ( .A1(instruction_1[21]), .A2(n8803), .ZN(n13843) );
  OAI22_X1 U17404 ( .A1(instruction_1[22]), .A2(n13843), .B1(n13843), .B2(
        n8806), .ZN(n13845) );
  XNOR2_X1 U17405 ( .A(rw_2[2]), .B(instruction_1[23]), .ZN(n13844) );
  NAND3_X1 U17406 ( .A1(n13846), .A2(n13845), .A3(n13844), .ZN(n13849) );
  XOR2_X1 U17407 ( .A(rw_2[3]), .B(instruction_1[24]), .Z(n13848) );
  XOR2_X1 U17408 ( .A(rw_2[4]), .B(instruction_1[25]), .Z(n13847) );
  NOR3_X1 U17409 ( .A1(n13849), .A2(n13848), .A3(n13847), .ZN(N19) );
  NOR2_X1 U17410 ( .A1(n8795), .A2(instruction_1[21]), .ZN(n13850) );
  OAI22_X1 U17411 ( .A1(n13850), .A2(n8805), .B1(rw_1[1]), .B2(n13850), .ZN(
        n13854) );
  AND2_X1 U17412 ( .A1(instruction_1[21]), .A2(n8795), .ZN(n13851) );
  OAI22_X1 U17413 ( .A1(instruction_1[22]), .A2(n13851), .B1(n13851), .B2(
        n8796), .ZN(n13853) );
  XNOR2_X1 U17414 ( .A(rw_1[2]), .B(instruction_1[23]), .ZN(n13852) );
  NAND3_X1 U17415 ( .A1(n13854), .A2(n13853), .A3(n13852), .ZN(n13857) );
  XOR2_X1 U17416 ( .A(rw_1[3]), .B(instruction_1[24]), .Z(n13856) );
  XOR2_X1 U17417 ( .A(rw_1[4]), .B(instruction_1[25]), .Z(n13855) );
  NOR3_X1 U17418 ( .A1(n13857), .A2(n13856), .A3(n13855), .ZN(N17) );
  INV_X4 U17419 ( .A(n382), .ZN(n16152) );
  INV_X4 U17420 ( .A(n380), .ZN(n16153) );
  INV_X4 U17421 ( .A(n378), .ZN(n16154) );
  INV_X4 U17422 ( .A(n376), .ZN(n16155) );
  INV_X4 U17423 ( .A(n374), .ZN(n16156) );
  INV_X4 U17424 ( .A(n372), .ZN(n16157) );
  INV_X4 U17425 ( .A(n366), .ZN(n16158) );
  INV_X4 U17426 ( .A(n364), .ZN(n16159) );
  INV_X4 U17427 ( .A(n362), .ZN(n16160) );
  INV_X4 U17428 ( .A(n360), .ZN(n16161) );
  INV_X4 U17429 ( .A(n358), .ZN(n16162) );
  INV_X4 U17430 ( .A(n356), .ZN(n16163) );
  INV_X4 U17431 ( .A(n354), .ZN(n16164) );
  INV_X4 U17432 ( .A(n352), .ZN(n16165) );
  INV_X4 U17433 ( .A(n350), .ZN(n16166) );
  INV_X4 U17434 ( .A(n348), .ZN(n16167) );
  INV_X4 U17435 ( .A(n346), .ZN(n16168) );
  INV_X4 U17436 ( .A(n344), .ZN(n16169) );
  INV_X4 U17437 ( .A(n342), .ZN(n16170) );
  INV_X4 U17438 ( .A(n340), .ZN(n16171) );
  INV_X4 U17439 ( .A(n338), .ZN(n16172) );
  INV_X4 U17440 ( .A(n330), .ZN(n16173) );
  INV_X4 U17441 ( .A(decode_N2), .ZN(n16174) );
  INV_X4 U17442 ( .A(decode_N4), .ZN(n16175) );
  INV_X4 U17443 ( .A(aluout_0[31]), .ZN(n16176) );
  INV_X4 U17444 ( .A(aluout_0[30]), .ZN(n16177) );
  INV_X4 U17445 ( .A(aluout_0[27]), .ZN(n16178) );
  INV_X4 U17446 ( .A(aluout_0[28]), .ZN(n16179) );
  INV_X4 U17447 ( .A(aluout_0[29]), .ZN(n16180) );
  INV_X4 U17448 ( .A(n3468), .ZN(n16181) );
  INV_X4 U17449 ( .A(n3472), .ZN(n16182) );
  INV_X4 U17450 ( .A(n2981), .ZN(n16183) );
  INV_X4 U17451 ( .A(n3482), .ZN(n16184) );
  INV_X4 U17452 ( .A(n3502), .ZN(n16185) );
  INV_X4 U17453 ( .A(n3509), .ZN(n16186) );
  INV_X4 U17454 ( .A(n3517), .ZN(n16187) );
  INV_X4 U17455 ( .A(n3523), .ZN(n16188) );
  INV_X4 U17456 ( .A(aluout_0[25]), .ZN(n16189) );
  INV_X4 U17457 ( .A(aluout_0[26]), .ZN(n16190) );
  INV_X4 U17458 ( .A(n3827), .ZN(n16191) );
  INV_X4 U17459 ( .A(n3974), .ZN(n16192) );
  INV_X4 U17460 ( .A(aluout_0[20]), .ZN(n16193) );
  INV_X4 U17461 ( .A(aluout_0[21]), .ZN(n16194) );
  INV_X4 U17462 ( .A(aluout_0[22]), .ZN(n16195) );
  INV_X4 U17463 ( .A(aluout_0[23]), .ZN(n16196) );
  INV_X4 U17464 ( .A(aluout_0[24]), .ZN(n16197) );
  INV_X4 U17465 ( .A(n4274), .ZN(n16198) );
  INV_X4 U17466 ( .A(n4280), .ZN(n16199) );
  INV_X4 U17467 ( .A(n4421), .ZN(n16200) );
  INV_X4 U17468 ( .A(n4554), .ZN(n16201) );
  INV_X4 U17469 ( .A(n4555), .ZN(n16202) );
  INV_X4 U17470 ( .A(n4286), .ZN(n16203) );
  INV_X4 U17471 ( .A(n4427), .ZN(n16204) );
  INV_X4 U17472 ( .A(n4561), .ZN(n16205) );
  INV_X4 U17473 ( .A(n4292), .ZN(n16206) );
  INV_X4 U17474 ( .A(n4433), .ZN(n16207) );
  INV_X4 U17475 ( .A(n4567), .ZN(n16208) );
  INV_X4 U17476 ( .A(aluout_0[19]), .ZN(n16209) );
  INV_X4 U17477 ( .A(aluout_0[18]), .ZN(n16210) );
  INV_X4 U17478 ( .A(aluout_0[17]), .ZN(n16211) );
  INV_X4 U17479 ( .A(aluout_0[0]), .ZN(n16212) );
  INV_X4 U17480 ( .A(n41), .ZN(n16213) );
  INV_X4 U17481 ( .A(N47), .ZN(n16214) );
  INV_X4 U17482 ( .A(n6186), .ZN(n16215) );
  INV_X4 U17483 ( .A(n6187), .ZN(n16216) );
  INV_X4 U17484 ( .A(fwdA[0]), .ZN(n16217) );
  INV_X4 U17485 ( .A(n20), .ZN(n16218) );
  INV_X4 U17486 ( .A(n19), .ZN(n16219) );
  INV_X4 U17487 ( .A(n18), .ZN(n16220) );
  INV_X4 U17488 ( .A(n17), .ZN(n16221) );
  INV_X4 U17489 ( .A(n16), .ZN(n16222) );
  INV_X4 U17490 ( .A(n15), .ZN(n16223) );
  INV_X4 U17491 ( .A(n34), .ZN(n16224) );
  INV_X4 U17492 ( .A(n35), .ZN(n16225) );
  INV_X4 U17493 ( .A(n36), .ZN(n16226) );
  INV_X4 U17494 ( .A(n37), .ZN(n16227) );
  INV_X4 U17495 ( .A(n30), .ZN(n16228) );
  INV_X4 U17496 ( .A(n31), .ZN(n16229) );
  INV_X4 U17497 ( .A(n32), .ZN(n16230) );
  INV_X4 U17498 ( .A(n33), .ZN(n16231) );
  INV_X4 U17499 ( .A(n26), .ZN(n16232) );
  INV_X4 U17500 ( .A(n27), .ZN(n16233) );
  INV_X4 U17501 ( .A(n28), .ZN(n16234) );
  INV_X4 U17502 ( .A(n29), .ZN(n16235) );
  INV_X4 U17503 ( .A(n22), .ZN(n16236) );
  INV_X4 U17504 ( .A(n23), .ZN(n16237) );
  INV_X4 U17505 ( .A(n24), .ZN(n16238) );
  INV_X4 U17506 ( .A(n25), .ZN(n16239) );
  INV_X4 U17507 ( .A(n45), .ZN(n16240) );
  INV_X4 U17508 ( .A(n44), .ZN(n16241) );
  INV_X4 U17509 ( .A(n42), .ZN(n16242) );
  INV_X4 U17510 ( .A(n43), .ZN(n16243) );
  INV_X4 U17511 ( .A(n38), .ZN(n16244) );
  INV_X4 U17512 ( .A(n39), .ZN(n16245) );
  INV_X4 U17513 ( .A(n40), .ZN(n16246) );
  INV_X4 U17514 ( .A(n49), .ZN(n16247) );
  INV_X4 U17515 ( .A(n48), .ZN(n16248) );
  INV_X4 U17516 ( .A(n47), .ZN(n16249) );
  INV_X4 U17517 ( .A(n46), .ZN(n16250) );
  INV_X4 U17518 ( .A(n53), .ZN(n16251) );
  INV_X4 U17519 ( .A(n52), .ZN(n16252) );
  INV_X4 U17520 ( .A(n51), .ZN(n16253) );
  INV_X4 U17521 ( .A(n50), .ZN(n16254) );
  INV_X4 U17522 ( .A(n2621), .ZN(n16255) );
  INV_X4 U17523 ( .A(aluout_0[9]), .ZN(n16256) );
  INV_X4 U17524 ( .A(n3294), .ZN(n16257) );
  INV_X4 U17525 ( .A(n3531), .ZN(n16258) );
  INV_X4 U17526 ( .A(n3537), .ZN(n16259) );
  INV_X4 U17527 ( .A(n3365), .ZN(n16260) );
  INV_X4 U17528 ( .A(n3300), .ZN(n16261) );
  INV_X4 U17529 ( .A(n3550), .ZN(n16262) );
  INV_X4 U17530 ( .A(n3357), .ZN(n16263) );
  INV_X4 U17531 ( .A(n3311), .ZN(n16264) );
  INV_X4 U17532 ( .A(n3870), .ZN(n16265) );
  INV_X4 U17533 ( .A(n4298), .ZN(n16266) );
  INV_X4 U17534 ( .A(n4304), .ZN(n16267) );
  INV_X4 U17535 ( .A(n4310), .ZN(n16268) );
  INV_X4 U17536 ( .A(n4171), .ZN(n16269) );
  INV_X4 U17537 ( .A(n4316), .ZN(n16270) );
  INV_X4 U17538 ( .A(n4036), .ZN(n16271) );
  INV_X4 U17539 ( .A(n4439), .ZN(n16272) );
  INV_X4 U17540 ( .A(n4573), .ZN(n16273) );
  INV_X4 U17541 ( .A(n4445), .ZN(n16274) );
  INV_X4 U17542 ( .A(n4579), .ZN(n16275) );
  INV_X4 U17543 ( .A(n4451), .ZN(n16276) );
  INV_X4 U17544 ( .A(n4585), .ZN(n16277) );
  INV_X4 U17545 ( .A(n4457), .ZN(n16278) );
  INV_X4 U17546 ( .A(n4591), .ZN(n16279) );
  INV_X4 U17547 ( .A(n4463), .ZN(n16280) );
  INV_X4 U17548 ( .A(n4597), .ZN(n16281) );
  INV_X4 U17549 ( .A(n4703), .ZN(n16282) );
  INV_X4 U17550 ( .A(n4825), .ZN(n16283) );
  INV_X4 U17551 ( .A(n4709), .ZN(n16284) );
  INV_X4 U17552 ( .A(n4831), .ZN(n16285) );
  INV_X4 U17553 ( .A(n4715), .ZN(n16286) );
  INV_X4 U17554 ( .A(n4837), .ZN(n16287) );
  INV_X4 U17555 ( .A(n4721), .ZN(n16288) );
  INV_X4 U17556 ( .A(n4843), .ZN(n16289) );
  INV_X4 U17557 ( .A(n4727), .ZN(n16290) );
  INV_X4 U17558 ( .A(n4849), .ZN(n16291) );
  INV_X4 U17559 ( .A(n4733), .ZN(n16292) );
  INV_X4 U17560 ( .A(n4855), .ZN(n16293) );
  INV_X4 U17561 ( .A(aluout_0[15]), .ZN(n16294) );
  INV_X4 U17562 ( .A(n5367), .ZN(n16295) );
  INV_X4 U17563 ( .A(aluout_0[16]), .ZN(n16296) );
  INV_X4 U17564 ( .A(n4975), .ZN(n16297) );
  INV_X4 U17565 ( .A(n5373), .ZN(n16298) );
  INV_X4 U17566 ( .A(n4981), .ZN(n16299) );
  INV_X4 U17567 ( .A(n5087), .ZN(n16300) );
  INV_X4 U17568 ( .A(n5188), .ZN(n16301) );
  INV_X4 U17569 ( .A(n5192), .ZN(n16302) );
  INV_X4 U17570 ( .A(n4987), .ZN(n16303) );
  INV_X4 U17571 ( .A(n5093), .ZN(n16304) );
  INV_X4 U17572 ( .A(n4993), .ZN(n16305) );
  INV_X4 U17573 ( .A(n5099), .ZN(n16306) );
  INV_X4 U17574 ( .A(n4999), .ZN(n16307) );
  INV_X4 U17575 ( .A(n5105), .ZN(n16308) );
  INV_X4 U17576 ( .A(n5205), .ZN(n16309) );
  INV_X4 U17577 ( .A(n5211), .ZN(n16310) );
  INV_X4 U17578 ( .A(aluout_0[12]), .ZN(n16311) );
  INV_X4 U17579 ( .A(aluout_0[14]), .ZN(n16312) );
  INV_X4 U17580 ( .A(aluout_0[13]), .ZN(n16313) );
  INV_X4 U17581 ( .A(n5545), .ZN(n16314) );
  INV_X4 U17582 ( .A(n5476), .ZN(n16315) );
  INV_X4 U17583 ( .A(aluout_0[11]), .ZN(n16316) );
  INV_X4 U17584 ( .A(n5726), .ZN(n16317) );
  INV_X4 U17585 ( .A(n5732), .ZN(n16318) );
  INV_X4 U17586 ( .A(aluout_0[10]), .ZN(n16319) );
  INV_X4 U17587 ( .A(n5730), .ZN(n16320) );
  INV_X4 U17588 ( .A(n2713), .ZN(n16321) );
  INV_X4 U17589 ( .A(n6076), .ZN(n16322) );
  INV_X4 U17590 ( .A(n5048), .ZN(n16323) );
  INV_X4 U17591 ( .A(aluout_0[8]), .ZN(n16324) );
  INV_X4 U17592 ( .A(n3353), .ZN(n16325) );
  INV_X4 U17593 ( .A(n5400), .ZN(n16326) );
  INV_X4 U17594 ( .A(n5482), .ZN(n16327) );
  INV_X4 U17595 ( .A(n5565), .ZN(n16328) );
  INV_X4 U17596 ( .A(n2760), .ZN(n16329) );
  INV_X4 U17597 ( .A(n5259), .ZN(n16330) );
  INV_X4 U17598 ( .A(n6025), .ZN(n16331) );
  INV_X4 U17599 ( .A(n5818), .ZN(n16332) );
  INV_X4 U17600 ( .A(aluout_0[5]), .ZN(n16333) );
  INV_X4 U17601 ( .A(n3313), .ZN(n16334) );
  INV_X4 U17602 ( .A(n3319), .ZN(n16335) );
  INV_X4 U17603 ( .A(n3349), .ZN(n16336) );
  INV_X4 U17604 ( .A(n3325), .ZN(n16337) );
  INV_X4 U17605 ( .A(n5344), .ZN(n16338) );
  INV_X4 U17606 ( .A(n5348), .ZN(n16339) );
  INV_X4 U17607 ( .A(n5571), .ZN(n16340) );
  INV_X4 U17608 ( .A(n5666), .ZN(n16341) );
  INV_X4 U17609 ( .A(n5744), .ZN(n16342) );
  INV_X4 U17610 ( .A(n5750), .ZN(n16343) );
  INV_X4 U17611 ( .A(n5845), .ZN(n16344) );
  INV_X4 U17612 ( .A(n5827), .ZN(n16345) );
  INV_X4 U17613 ( .A(n5843), .ZN(n16346) );
  INV_X4 U17614 ( .A(n2740), .ZN(n16347) );
  INV_X4 U17615 ( .A(n5858), .ZN(n16348) );
  INV_X4 U17616 ( .A(aluout_0[7]), .ZN(n16349) );
  INV_X4 U17617 ( .A(n2767), .ZN(n16350) );
  INV_X4 U17618 ( .A(n5854), .ZN(n16351) );
  INV_X4 U17619 ( .A(aluout_0[6]), .ZN(n16352) );
  INV_X4 U17620 ( .A(n2797), .ZN(n16353) );
  INV_X4 U17621 ( .A(n2840), .ZN(n16354) );
  INV_X4 U17622 ( .A(n5778), .ZN(n16355) );
  INV_X4 U17623 ( .A(n2813), .ZN(n16356) );
  INV_X4 U17624 ( .A(n267), .ZN(n16357) );
  INV_X4 U17625 ( .A(n3196), .ZN(n16358) );
  INV_X4 U17626 ( .A(n6069), .ZN(n16359) );
  INV_X4 U17627 ( .A(n5451), .ZN(n16360) );
  INV_X4 U17628 ( .A(n3625), .ZN(n16361) );
  INV_X4 U17629 ( .A(n5535), .ZN(n16362) );
  INV_X4 U17630 ( .A(n3939), .ZN(n16363) );
  INV_X4 U17631 ( .A(n6070), .ZN(n16364) );
  INV_X4 U17632 ( .A(n5633), .ZN(n16365) );
  INV_X4 U17633 ( .A(n4237), .ZN(n16366) );
  INV_X4 U17634 ( .A(n5717), .ZN(n16367) );
  INV_X4 U17635 ( .A(n5795), .ZN(n16368) );
  INV_X4 U17636 ( .A(n4522), .ZN(n16369) );
  INV_X4 U17637 ( .A(n5780), .ZN(n16370) );
  INV_X4 U17638 ( .A(stallack), .ZN(n16371) );
  INV_X4 U17639 ( .A(n3345), .ZN(n16372) );
  INV_X4 U17640 ( .A(n3920), .ZN(n16373) );
  INV_X4 U17641 ( .A(n4073), .ZN(n16374) );
  INV_X4 U17642 ( .A(n3595), .ZN(n16375) );
  INV_X4 U17643 ( .A(n3599), .ZN(n16376) );
  INV_X4 U17644 ( .A(n4209), .ZN(n16377) );
  INV_X4 U17645 ( .A(n4755), .ZN(n16378) );
  INV_X4 U17646 ( .A(n3585), .ZN(n16379) );
  INV_X4 U17647 ( .A(n3589), .ZN(n16380) );
  INV_X4 U17648 ( .A(n4197), .ZN(n16381) );
  INV_X4 U17649 ( .A(n4201), .ZN(n16382) );
  INV_X4 U17650 ( .A(n3438), .ZN(n16383) );
  INV_X4 U17651 ( .A(n2906), .ZN(n16384) );
  INV_X4 U17652 ( .A(n2912), .ZN(n16385) );
  INV_X4 U17653 ( .A(n5787), .ZN(n16386) );
  INV_X4 U17654 ( .A(aluout_0[3]), .ZN(n16387) );
  INV_X4 U17655 ( .A(n6103), .ZN(n16388) );
  INV_X4 U17656 ( .A(n4756), .ZN(n16389) );
  INV_X4 U17657 ( .A(n4627), .ZN(n16390) );
  INV_X4 U17658 ( .A(n4057), .ZN(n16391) );
  INV_X4 U17659 ( .A(n3762), .ZN(n16392) );
  INV_X4 U17660 ( .A(n4063), .ZN(n16393) );
  INV_X4 U17661 ( .A(n4355), .ZN(n16394) );
  INV_X4 U17662 ( .A(n4633), .ZN(n16395) );
  INV_X4 U17663 ( .A(n5614), .ZN(n16396) );
  INV_X4 U17664 ( .A(aluout_0[1]), .ZN(n16397) );
  INV_X4 U17665 ( .A(n4943), .ZN(n16398) );
  INV_X4 U17666 ( .A(n5528), .ZN(n16399) );
  INV_X4 U17667 ( .A(aluout_0[2]), .ZN(n16400) );
  INV_X4 U17668 ( .A(n5359), .ZN(n16401) );
  INV_X4 U17669 ( .A(n5650), .ZN(n16402) );
  INV_X4 U17670 ( .A(aluout_0[4]), .ZN(n16403) );
  INV_X4 U17671 ( .A(n4884), .ZN(n16404) );
  INV_X4 U17672 ( .A(n4760), .ZN(n16405) );
  INV_X4 U17673 ( .A(n4803), .ZN(n16407) );
  INV_X4 U17674 ( .A(n4917), .ZN(n16408) );
  INV_X4 U17675 ( .A(n4537), .ZN(n16410) );
  INV_X4 U17676 ( .A(n4673), .ZN(n16411) );
  INV_X4 U17677 ( .A(n5062), .ZN(n16412) );
  INV_X4 U17678 ( .A(n2817), .ZN(n16413) );
  INV_X4 U17679 ( .A(n5606), .ZN(n16414) );
  INV_X4 U17680 ( .A(n5440), .ZN(n16415) );
  INV_X4 U17681 ( .A(n5800), .ZN(n16416) );
  INV_X4 U17682 ( .A(n4790), .ZN(n16417) );
  INV_X4 U17683 ( .A(n5272), .ZN(n16418) );
  INV_X4 U17684 ( .A(n5360), .ZN(n16419) );
  INV_X4 U17685 ( .A(n3442), .ZN(n16420) );
  INV_X4 U17686 ( .A(n6160), .ZN(n16421) );
  INV_X4 U17687 ( .A(n6073), .ZN(n16422) );
  INV_X4 U17688 ( .A(n6085), .ZN(n16423) );
  INV_X4 U17689 ( .A(n2970), .ZN(n16424) );
  INV_X4 U17690 ( .A(n3451), .ZN(n16425) );
  INV_X4 U17691 ( .A(n3455), .ZN(n16426) );
  INV_X4 U17692 ( .A(n3209), .ZN(n16427) );
  INV_X4 U17693 ( .A(n3952), .ZN(n16428) );
  INV_X4 U17694 ( .A(n2946), .ZN(n16429) );
  INV_X4 U17695 ( .A(n4533), .ZN(n16430) );
  INV_X4 U17696 ( .A(n4252), .ZN(n16432) );
  INV_X4 U17697 ( .A(n4248), .ZN(n16434) );
  INV_X4 U17698 ( .A(n3227), .ZN(n16436) );
  INV_X4 U17699 ( .A(n6128), .ZN(n16437) );
  INV_X4 U17700 ( .A(n6078), .ZN(n16438) );
  INV_X4 U17701 ( .A(n4114), .ZN(n16439) );
  INV_X4 U17702 ( .A(n4259), .ZN(n16440) );
  INV_X4 U17703 ( .A(n4794), .ZN(n16441) );
  INV_X4 U17704 ( .A(n4662), .ZN(n16442) );
  INV_X4 U17705 ( .A(n4526), .ZN(n16443) );
  INV_X4 U17706 ( .A(n3426), .ZN(n16444) );
  INV_X4 U17707 ( .A(n3802), .ZN(n16445) );
  INV_X4 U17708 ( .A(n3651), .ZN(n16446) );
  INV_X4 U17709 ( .A(n2823), .ZN(n16447) );
  INV_X4 U17710 ( .A(n6032), .ZN(n16450) );
  INV_X4 U17711 ( .A(n2861), .ZN(n16451) );
  INV_X4 U17712 ( .A(n3231), .ZN(n16452) );
  INV_X4 U17713 ( .A(n3964), .ZN(n16453) );
  INV_X4 U17714 ( .A(n5708), .ZN(n16454) );
  INV_X4 U17715 ( .A(n5641), .ZN(n16457) );
  INV_X4 U17716 ( .A(n4955), .ZN(n16459) );
  INV_X4 U17717 ( .A(n5934), .ZN(n16460) );
  INV_X4 U17718 ( .A(n6014), .ZN(n16461) );
  INV_X4 U17719 ( .A(n4245), .ZN(n16462) );
  INV_X4 U17720 ( .A(n2894), .ZN(n16463) );
  INV_X4 U17721 ( .A(n3404), .ZN(n16464) );
  INV_X4 U17722 ( .A(n4386), .ZN(n16465) );
  INV_X4 U17723 ( .A(n2856), .ZN(n16466) );
  INV_X4 U17724 ( .A(n3234), .ZN(n16467) );
  INV_X4 U17725 ( .A(n4666), .ZN(n16468) );
  INV_X4 U17726 ( .A(n2706), .ZN(n16470) );
  INV_X4 U17727 ( .A(n5229), .ZN(n16472) );
  INV_X4 U17728 ( .A(n5230), .ZN(n16473) );
  INV_X4 U17729 ( .A(n2851), .ZN(n16474) );
  INV_X4 U17730 ( .A(n5683), .ZN(n16475) );
  INV_X4 U17731 ( .A(n5687), .ZN(n16476) );
  INV_X4 U17732 ( .A(n5893), .ZN(n16477) );
  INV_X4 U17733 ( .A(n6124), .ZN(n16478) );
  INV_X4 U17734 ( .A(n6034), .ZN(n16479) );
  INV_X4 U17735 ( .A(n3335), .ZN(n16480) );
  INV_X4 U17736 ( .A(n3336), .ZN(n16481) );
  INV_X4 U17737 ( .A(n5052), .ZN(n16482) );
  INV_X4 U17738 ( .A(n5026), .ZN(n16483) );
  INV_X4 U17739 ( .A(n5418), .ZN(n16484) );
  INV_X4 U17740 ( .A(n5238), .ZN(n16485) );
  INV_X4 U17741 ( .A(n3965), .ZN(n16486) );
  INV_X4 U17742 ( .A(n5587), .ZN(n16487) );
  INV_X4 U17743 ( .A(n4941), .ZN(n16488) );
  INV_X4 U17744 ( .A(n2839), .ZN(n16489) );
  INV_X4 U17745 ( .A(n5174), .ZN(n16490) );
  INV_X4 U17746 ( .A(n4683), .ZN(n16491) );
  INV_X4 U17747 ( .A(n4246), .ZN(n16492) );
  INV_X4 U17748 ( .A(n3643), .ZN(n16493) );
  INV_X4 U17749 ( .A(n3803), .ZN(n16494) );
  INV_X4 U17750 ( .A(n2790), .ZN(n16495) );
  INV_X4 U17751 ( .A(n4405), .ZN(n16496) );
  INV_X4 U17752 ( .A(n5899), .ZN(n16497) );
  INV_X4 U17753 ( .A(n5917), .ZN(n16498) );
  INV_X4 U17754 ( .A(n5970), .ZN(n16499) );
  INV_X4 U17755 ( .A(n5983), .ZN(n16500) );
  INV_X4 U17756 ( .A(n5995), .ZN(n16501) );
  INV_X4 U17757 ( .A(n4390), .ZN(n16502) );
  INV_X4 U17758 ( .A(n5071), .ZN(n16503) );
  INV_X4 U17759 ( .A(n6010), .ZN(n16504) );
  INV_X4 U17760 ( .A(n4101), .ZN(n16505) );
  INV_X4 U17761 ( .A(n3652), .ZN(n16506) );
  INV_X4 U17762 ( .A(n4261), .ZN(n16507) );
  INV_X4 U17763 ( .A(n3242), .ZN(n16508) );
  INV_X4 U17764 ( .A(n2784), .ZN(n16509) );
  INV_X4 U17765 ( .A(n3241), .ZN(n16510) );
  INV_X4 U17766 ( .A(n3640), .ZN(n16511) );
  INV_X4 U17767 ( .A(n5643), .ZN(n16512) );
  INV_X4 U17768 ( .A(n3420), .ZN(n16513) );
  INV_X4 U17769 ( .A(n2816), .ZN(n16514) );
  INV_X4 U17770 ( .A(n3445), .ZN(n16515) );
  INV_X4 U17771 ( .A(n6020), .ZN(n16516) );
  INV_X4 U17772 ( .A(n3443), .ZN(n16517) );
  INV_X4 U17773 ( .A(n4530), .ZN(n16518) );
  INV_X4 U17774 ( .A(n3245), .ZN(n16519) );
  INV_X4 U17775 ( .A(n3247), .ZN(n16520) );
  INV_X4 U17776 ( .A(n5262), .ZN(n16521) );
  INV_X4 U17777 ( .A(n5590), .ZN(n16522) );
  INV_X4 U17778 ( .A(n5421), .ZN(n16523) );
  INV_X4 U17779 ( .A(n2917), .ZN(n16524) );
  INV_X4 U17780 ( .A(n4766), .ZN(n16525) );
  INV_X4 U17781 ( .A(n4492), .ZN(n16526) );
  INV_X4 U17782 ( .A(n4206), .ZN(n16527) );
  INV_X4 U17783 ( .A(n3908), .ZN(n16528) );
  INV_X4 U17784 ( .A(n2884), .ZN(n16529) );
  INV_X4 U17785 ( .A(n2880), .ZN(n16530) );
  INV_X4 U17786 ( .A(n2882), .ZN(n16531) );
  INV_X4 U17787 ( .A(n2885), .ZN(n16532) );
  INV_X4 U17788 ( .A(n6044), .ZN(n16533) );
  INV_X4 U17789 ( .A(n4490), .ZN(n16534) );
  INV_X4 U17790 ( .A(n4764), .ZN(n16535) );
  INV_X4 U17791 ( .A(n5131), .ZN(n16536) );
  INV_X4 U17792 ( .A(n3641), .ZN(n16537) );
  INV_X4 U17793 ( .A(n4205), .ZN(n16538) );
  INV_X4 U17794 ( .A(n3408), .ZN(n16539) );
  INV_X4 U17795 ( .A(n3412), .ZN(n16540) );
  INV_X4 U17796 ( .A(n3411), .ZN(n16541) );
  INV_X4 U17797 ( .A(n5692), .ZN(n16542) );
  INV_X4 U17798 ( .A(n5505), .ZN(n16543) );
  INV_X4 U17799 ( .A(n5326), .ZN(n16544) );
  INV_X4 U17800 ( .A(n5646), .ZN(n16545) );
  INV_X4 U17801 ( .A(n5616), .ZN(n16546) );
  INV_X4 U17802 ( .A(fwdB[1]), .ZN(n16547) );
  INV_X4 U17803 ( .A(n3429), .ZN(n16549) );
  INV_X4 U17804 ( .A(n21), .ZN(n16550) );
  INV_X4 U17805 ( .A(n3403), .ZN(n16551) );
  INV_X4 U17806 ( .A(n2578), .ZN(n16552) );
  INV_X4 U17807 ( .A(n2581), .ZN(n16553) );
  INV_X4 U17808 ( .A(n2583), .ZN(n16554) );
  INV_X4 U17809 ( .A(n2585), .ZN(n16555) );
  INV_X4 U17810 ( .A(n2587), .ZN(n16556) );
  INV_X4 U17811 ( .A(n2589), .ZN(n16557) );
  INV_X4 U17812 ( .A(n2591), .ZN(n16558) );
  INV_X4 U17813 ( .A(n2593), .ZN(n16559) );
  INV_X4 U17814 ( .A(n2595), .ZN(n16560) );
  INV_X4 U17815 ( .A(n2597), .ZN(n16561) );
  INV_X4 U17816 ( .A(n2599), .ZN(n16562) );
  INV_X4 U17817 ( .A(n2601), .ZN(n16563) );
  INV_X4 U17818 ( .A(n2603), .ZN(n16564) );
  INV_X4 U17819 ( .A(n2605), .ZN(n16565) );
  INV_X4 U17820 ( .A(n2607), .ZN(n16566) );
  INV_X4 U17821 ( .A(n2609), .ZN(n16567) );
  INV_X4 U17822 ( .A(n2611), .ZN(n16568) );
  INV_X4 U17823 ( .A(n2613), .ZN(n16569) );
  INV_X4 U17824 ( .A(n2615), .ZN(n16570) );
  INV_X4 U17825 ( .A(n2617), .ZN(n16571) );
  INV_X4 U17826 ( .A(n2619), .ZN(n16572) );
  INV_X4 U17827 ( .A(n2623), .ZN(n16573) );
  INV_X4 U17828 ( .A(n2625), .ZN(n16574) );
  INV_X4 U17829 ( .A(n2627), .ZN(n16575) );
  INV_X4 U17830 ( .A(n2629), .ZN(n16576) );
  INV_X4 U17831 ( .A(n2631), .ZN(n16577) );
  INV_X4 U17832 ( .A(n2633), .ZN(n16578) );
  INV_X4 U17833 ( .A(n2635), .ZN(n16579) );
  INV_X4 U17834 ( .A(n2637), .ZN(n16580) );
  INV_X4 U17835 ( .A(n2639), .ZN(n16581) );
  INV_X4 U17836 ( .A(n2641), .ZN(n16582) );
  INV_X4 U17837 ( .A(n2654), .ZN(n16583) );
  INV_X4 U17838 ( .A(n2662), .ZN(n16584) );
  INV_X4 U17839 ( .A(n2663), .ZN(n16585) );
  INV_X4 U17840 ( .A(n2647), .ZN(n16586) );
  INV_X4 U17841 ( .A(n2675), .ZN(n16587) );
  INV_X4 U17842 ( .A(n138), .ZN(n16588) );
  INV_X4 U17843 ( .A(n283), .ZN(n16589) );
  INV_X4 U17844 ( .A(n145), .ZN(n16590) );
  INV_X4 U17845 ( .A(n305), .ZN(n16591) );
  INV_X4 U17846 ( .A(n293), .ZN(n16592) );
  INV_X4 U17847 ( .A(n2660), .ZN(n16593) );
  INV_X4 U17848 ( .A(n161), .ZN(n16594) );
  INV_X4 U17849 ( .A(n2692), .ZN(n16595) );
  INV_X4 U17850 ( .A(n2690), .ZN(n16596) );
  INV_X4 U17851 ( .A(n292), .ZN(n16597) );
  INV_X4 U17852 ( .A(n160), .ZN(n16598) );
  INV_X4 U17853 ( .A(n2689), .ZN(n16599) );
  INV_X4 U17854 ( .A(n306), .ZN(n16600) );
  INV_X4 U17855 ( .A(n2644), .ZN(n16601) );
  INV_X4 U17856 ( .A(n149), .ZN(n16602) );
  INV_X4 U17857 ( .A(n2695), .ZN(n16603) );
  INV_X4 U17858 ( .A(n2688), .ZN(n16604) );
  INV_X4 U17859 ( .A(n2691), .ZN(n16605) );
endmodule

